`define UNIT_DELAY #1
`define USE_POWER_PINS
`define FUNCTIONAL
`include "libs.ref/sky130_fd_sc_hd/verilog/primitives.v"
`include "libs.ref/sky130_fd_sc_hd/verilog/sky130_fd_sc_hd.v"

module fib (clk,
    rdy_in,
    rdy_out,
    rst_n,
    vld_in,
    vld_out,
    VPWR,
    VGND,
    fib_in,
    fib_out);
 input clk;
 output rdy_in;
 input rdy_out;
 input rst_n;
 input vld_in;
 output vld_out;
 inout VPWR;
 inout VGND;
 input [7:0] fib_in;
 output [31:0] fib_out;

 wire fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D;
 wire fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1;
 wire \iters[0] ;
 wire \iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \iters[1] ;
 wire \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \iters[2] ;
 wire \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \iters[3] ;
 wire \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ;
 wire \iters[4] ;
 wire \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \iters[5] ;
 wire \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \iters[6] ;
 wire \iters[6]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \iters[6]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ;
 wire \iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[7] ;
 wire \iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \iters[7]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \iters[7]_sky130_fd_sc_hd__o21a_2_B1_A2 ;
 wire \iters[7]_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \prev1[0] ;
 wire \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev1[10] ;
 wire \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \prev1[11] ;
 wire \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[12] ;
 wire \prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[13] ;
 wire \prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[14] ;
 wire \prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[15] ;
 wire \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X_A1 ;
 wire \prev1[16] ;
 wire \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[17] ;
 wire \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[18] ;
 wire \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ;
 wire \prev1[19] ;
 wire \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[1] ;
 wire \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[20] ;
 wire \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ;
 wire \prev1[21] ;
 wire \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[22] ;
 wire \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[23] ;
 wire \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[24] ;
 wire \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[25] ;
 wire \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X_A2 ;
 wire \prev1[26] ;
 wire \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[27] ;
 wire \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[28] ;
 wire \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ;
 wire \prev1[29] ;
 wire \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[2] ;
 wire \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[30] ;
 wire \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X_A ;
 wire \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[31] ;
 wire \prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[3] ;
 wire \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[4] ;
 wire \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ;
 wire \prev1[5] ;
 wire \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[6] ;
 wire \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[7] ;
 wire \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev1[8] ;
 wire \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A ;
 wire \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X_B ;
 wire \prev1[9] ;
 wire \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ;
 wire \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \prev2[0] ;
 wire \prev2[0]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[0]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[10] ;
 wire \prev2[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[10]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \prev2[11] ;
 wire \prev2[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X ;
 wire \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X_sky130_fd_sc_hd__and3b_2_B_X ;
 wire \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \prev2[12] ;
 wire \prev2[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_A3 ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_B1 ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_C1 ;
 wire \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_X ;
 wire \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ;
 wire \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D ;
 wire \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ;
 wire \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or3_2_C_X ;
 wire \prev2[13] ;
 wire \prev2[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[13]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \prev2[14] ;
 wire \prev2[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[15] ;
 wire \prev2[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[16] ;
 wire \prev2[16]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \prev2[17] ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_B1 ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_A2 ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1 ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \prev2[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1 ;
 wire \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \prev2[18] ;
 wire \prev2[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[18]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[19] ;
 wire \prev2[19]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[1] ;
 wire \prev2[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[1]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[1]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ;
 wire \prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \prev2[20] ;
 wire \prev2[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[20]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \prev2[21] ;
 wire \prev2[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_C ;
 wire \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_X ;
 wire \prev2[22] ;
 wire \prev2[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[22]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \prev2[23] ;
 wire \prev2[23]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[24] ;
 wire \prev2[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[25] ;
 wire \prev2[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_B ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ;
 wire \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \prev2[26] ;
 wire \prev2[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[26]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[27] ;
 wire \prev2[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_B1 ;
 wire \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ;
 wire \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A ;
 wire \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[28] ;
 wire \prev2[28]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ;
 wire \prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \prev2[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[29] ;
 wire \prev2[29]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[29]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ;
 wire \prev2[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[2] ;
 wire \prev2[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[2]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[30] ;
 wire \prev2[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[30]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[30]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[30]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \prev2[31] ;
 wire \prev2[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \prev2[3] ;
 wire \prev2[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X ;
 wire \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ;
 wire \prev2[3]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[4] ;
 wire \prev2[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[4]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[5] ;
 wire \prev2[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ;
 wire \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1 ;
 wire \prev2[6] ;
 wire \prev2[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[6]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \prev2[7] ;
 wire \prev2[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[7]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[8] ;
 wire \prev2[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[8]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \prev2[9] ;
 wire \prev2[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \prev2[9]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire rdy_in_sky130_fd_sc_hd__dfstp_2_Q_D;
 wire rdy_out_sky130_fd_sc_hd__o21ai_2_A2_B1;
 wire \state[2] ;
 wire \state[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ;
 wire \state[2]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \state[2]_sky130_fd_sc_hd__o211ai_2_A1_Y ;
 wire \state[2]_sky130_fd_sc_hd__o21a_2_B1_A1 ;
 wire \state[2]_sky130_fd_sc_hd__o21a_2_B1_A2 ;
 wire \state[2]_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \target_iters[0] ;
 wire \target_iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[1] ;
 wire \target_iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[1]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[2] ;
 wire \target_iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[2]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[3] ;
 wire \target_iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[3]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[4] ;
 wire \target_iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[4]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[5] ;
 wire \target_iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[5]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[6] ;
 wire \target_iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[6]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \target_iters[7] ;
 wire \target_iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \target_iters[7]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire vld_in_sky130_fd_sc_hd__and3_2_B_X;
 wire vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y;
 wire vld_out_sky130_fd_sc_hd__dfrtp_2_Q_D;
 wire vld_out_sky130_fd_sc_hd__inv_2_A_Y;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net85;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net84;
 wire net86;
 wire net100;
 wire net101;
 wire net103;

 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X (.A(\prev1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_1 (.A(\prev1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_10 (.A(\prev1[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_11 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_12 (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_13 (.A(\prev1[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_14 (.A(\prev1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_15 (.A(\prev1[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_16 (.A(\prev1[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_17 (.A(\prev1[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_18 (.A(\prev1[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_19 (.A(\prev1[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_2 (.A(\prev1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_20 (.A(\prev1[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_21 (.A(\prev1[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_22 (.A(\prev1[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_23 (.A(\prev1[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_24 (.A(\prev1[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_25 (.A(\prev1[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_26 (.A(\prev1[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_27 (.A(\prev1[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_28 (.A(\prev1[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_29 (.A(\prev1[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_3 (.A(\prev1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_30 (.A(\prev1[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_4 (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_5 (.A(\prev1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_6 (.A(\prev1[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_7 (.A(\prev1[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_8 (.A(\prev1[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 fib_out_sky130_fd_sc_hd__buf_2_X_9 (.A(\prev1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__dfrtp_1 fib_out_sky130_fd_sc_hd__dfrtp_2_Q (.CLK(clknet_3_6__leaf_clk),
    .D(fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net12));
 sky130_fd_sc_hd__a22o_1 fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X (.A1(net120),
    .A2(net60),
    .B1(fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D));
 sky130_fd_sc_hd__dfxtp_2 \iters[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[0] ));
 sky130_fd_sc_hd__inv_2 \iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__inv_2_Y  (.A(\iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__inv_2_Y_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__mux2_1_X  (.A0(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .S(\iters[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__dfxtp_1 \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[1] ));
 sky130_fd_sc_hd__a32o_1 \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A2(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(\iters[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or2_2_X  (.A(\iters[0] ),
    .B(\iters[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand2_1 \iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nand2_2_Y  (.A(\iters[0] ),
    .B(\iters[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfxtp_2 \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[2] ));
 sky130_fd_sc_hd__a32o_1 \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A2(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(\iters[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\iters[0] ),
    .B(\iters[1] ),
    .C(\iters[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\iters[0] ),
    .A2(\iters[1] ),
    .B1(\iters[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfxtp_1 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[3] ));
 sky130_fd_sc_hd__a32o_1 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A2(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a31o_2_X  (.A1(\iters[0] ),
    .A2(\iters[1] ),
    .A3(\iters[2] ),
    .B1(\iters[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__inv_2 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y  (.A(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__and2_1 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B  (.A(\iters[4] ),
    .B(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and4_1 \iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and4_2_X  (.A(\iters[0] ),
    .B(\iters[1] ),
    .C(\iters[2] ),
    .D(\iters[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__dfxtp_1 \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[4] ));
 sky130_fd_sc_hd__a32o_1 \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A2(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or2_2_X  (.A(\iters[4] ),
    .B(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__inv_2 \iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y  (.A(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfxtp_1 \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[5] ));
 sky130_fd_sc_hd__a32o_1 \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A2(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or2_2_X  (.A(\iters[5] ),
    .B(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand2_1 \iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nand2_2_Y  (.A(\iters[5] ),
    .B(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__a31o_1 \iters[6]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\iters[5] ),
    .A2(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A3(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\iters[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[6]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \iters[6]_sky130_fd_sc_hd__and3_2_B  (.A(\iters[5] ),
    .B(\iters[6] ),
    .C(\iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[6]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .B(\iters[6]_sky130_fd_sc_hd__and3_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[7]_sky130_fd_sc_hd__o21a_2_B1_A2 ));
 sky130_fd_sc_hd__inv_2 \iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__inv_2_Y  (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__dfxtp_1 \iters[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[6] ));
 sky130_fd_sc_hd__o21a_1 \iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\iters[7]_sky130_fd_sc_hd__o21a_2_B1_A2 ),
    .B1(\iters[6]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \iters[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\iters[7] ));
 sky130_fd_sc_hd__a31o_1 \iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X  (.A1(\iters[7]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .A3(\iters[6]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\iters[7]_sky130_fd_sc_hd__o21a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \iters[7]_sky130_fd_sc_hd__inv_2_A  (.A(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\iters[7]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \iters[7]_sky130_fd_sc_hd__o21a_2_B1  (.A1(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\iters[7]_sky130_fd_sc_hd__o21a_2_B1_A2 ),
    .B1(\iters[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\iters[7]_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[0] ));
 sky130_fd_sc_hd__o22a_1 \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X  (.A1(net166),
    .A2(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__inv_2_Y  (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nand2_2 \prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B  (.A(net69),
    .B(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[0]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[10] ));
 sky130_fd_sc_hd__a32o_1 \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net50),
    .A2(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1(net59),
    .B2(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .A2(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X_B ),
    .B1(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[11] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[11] ),
    .B2(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X  (.A1(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A3(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[11]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[12] ));
 sky130_fd_sc_hd__a32o_1 \prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net52),
    .A2(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net60),
    .B2(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[13] ));
 sky130_fd_sc_hd__a32o_1 \prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net49),
    .A2(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net57),
    .B2(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_2 \prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[14] ));
 sky130_fd_sc_hd__a32o_1 \prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net49),
    .A2(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net57),
    .B2(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[15] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[15] ),
    .B2(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X_A1 ),
    .A2(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X  (.A1(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X_A1 ),
    .A2(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(net100),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__nand2_1 \prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X_A1_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev1[14] ),
    .B(\prev2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X_A1 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[16] ));
 sky130_fd_sc_hd__a32o_1 \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net50),
    .A2(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net59),
    .B2(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or2_2_X  (.A(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1 ),
    .B(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand2_1 \prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1 ),
    .B(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[16]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[17] ));
 sky130_fd_sc_hd__a32o_1 \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net47),
    .A2(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net55),
    .B2(\prev1[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_B1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[18] ));
 sky130_fd_sc_hd__a32o_1 \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net47),
    .A2(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net55),
    .B2(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__or2_4 \prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X  (.A(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[19] ));
 sky130_fd_sc_hd__a32o_1 \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net46),
    .A2(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net54),
    .B2(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__o211ai_1 \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__o211ai_2_Y  (.A1(\prev2[19]_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C1(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a211o_2_X  (.A1(\prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[19]_sky130_fd_sc_hd__and2_2_B_X ),
    .C1(\prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[19]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[1] ));
 sky130_fd_sc_hd__a32o_1 \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net52),
    .A2(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net60),
    .B2(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__inv_2_Y  (.A(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[20] ));
 sky130_fd_sc_hd__a22o_1 \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\prev1[20] ),
    .A2(net55),
    .B1(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1 ),
    .A2(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a31oi_1 \prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2_sky130_fd_sc_hd__a31oi_2_Y  (.A1(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1 ),
    .A3(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[21] ));
 sky130_fd_sc_hd__a32o_1 \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net46),
    .A2(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net54),
    .B2(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B1(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand3_1 \prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .C(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[22] ));
 sky130_fd_sc_hd__a32o_1 \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net46),
    .A2(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net54),
    .B2(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .C(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[21]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .B1(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[23] ));
 sky130_fd_sc_hd__a32o_1 \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net46),
    .A2(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net54),
    .B2(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__o211ai_1 \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__o211ai_2_Y  (.A1(\prev2[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C1(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a211o_2_X  (.A1(\prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[22]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .C1(\prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[23]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[24] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[24] ),
    .B2(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .B(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__nand2_1 \prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__nand2_2_Y  (.A(net46),
    .B(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X_A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[25] ));
 sky130_fd_sc_hd__a32o_1 \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net48),
    .A2(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net56),
    .B2(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\prev1[24] ),
    .A2(\prev2[24] ),
    .B1(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .B2(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ),
    .C1(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21bo_1 \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X  (.A1(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N ),
    .A2(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X_A2 ),
    .B1_N(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__nand2_1 \prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X_A2_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .B(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21bo_2_X_A2 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[26] ));
 sky130_fd_sc_hd__a32o_1 \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net48),
    .A2(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net56),
    .B2(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .C(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[25]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[27] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[27] ),
    .B2(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X  (.A1(\prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[26]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[27]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[28] ));
 sky130_fd_sc_hd__a22o_1 \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(net188),
    .A2(net56),
    .B1(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ),
    .B(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__o21a_1 \prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2_sky130_fd_sc_hd__o21a_2_X  (.A1(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ),
    .A2(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[28]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[29] ));
 sky130_fd_sc_hd__a32o_1 \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net48),
    .A2(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net56),
    .B2(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[2] ));
 sky130_fd_sc_hd__a32o_1 \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net50),
    .A2(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or2_2_X  (.A(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .B(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand2_1 \prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .B(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[30] ));
 sky130_fd_sc_hd__a32o_1 \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net48),
    .A2(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .B1(net56),
    .B2(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__or3_1 \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X  (.A(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\prev2[30]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__o21ai_4 \prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X_A ),
    .A2(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\prev2[30]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[31] ));
 sky130_fd_sc_hd__a2bb2o_4 \prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .A2_N(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .B1(\prev1[31] ),
    .B2(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[3] ));
 sky130_fd_sc_hd__a32o_1 \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net50),
    .A2(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .C(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[2]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .B1(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[3]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[4] ));
 sky130_fd_sc_hd__a32o_1 \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net51),
    .A2(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__or2_1 \prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X  (.A(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[5] ));
 sky130_fd_sc_hd__a32o_1 \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net51),
    .A2(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .C(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[6] ));
 sky130_fd_sc_hd__a32o_1 \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net51),
    .A2(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand3_1 \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y  (.A(\prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .C(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[5]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[7] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[7] ),
    .B2(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X  (.A1(\prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[6]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[8] ));
 sky130_fd_sc_hd__a32o_1 \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X  (.A1(net51),
    .A2(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net58),
    .B2(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__or2_1 \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X  (.A(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__and2_1 \prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X  (.A(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .B(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__dfrtp_1 \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev1[9] ));
 sky130_fd_sc_hd__a2bb2o_1 \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ),
    .A2_N(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\prev1[9] ),
    .B2(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__a31o_2_X  (.A1(\prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[9]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a22o_1 \prev2[0]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[0] ),
    .A2(net52),
    .B1(net60),
    .B2(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_4 \prev2[0]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[0] ),
    .B(\prev2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[0]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[0]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(net150),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[0] ));
 sky130_fd_sc_hd__nor2_1 \prev2[0]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[0] ),
    .B(\prev2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[0]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[0]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\prev2[0]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[0]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(fib_out_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1));
 sky130_fd_sc_hd__a22o_1 \prev2[10]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net190),
    .A2(net50),
    .B1(net59),
    .B2(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[10]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev2[10]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[10] ));
 sky130_fd_sc_hd__nand2_1 \prev2[10]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[10] ),
    .B(\prev2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[10]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[10] ),
    .B(\prev2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\prev1[10]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__nand3_2_Y_A ),
    .A2(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .B1(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[11]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[11] ),
    .A2(net52),
    .B1(net60),
    .B2(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[11]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev2[11]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[11] ));
 sky130_fd_sc_hd__nand2_1 \prev2[11]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[11] ),
    .B(\prev2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_1 \prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[11]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[11] ),
    .B(\prev2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a211o_1 \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1  (.A1(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ),
    .C1(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X ));
 sky130_fd_sc_hd__and3b_1 \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X_sky130_fd_sc_hd__and3b_2_B  (.A_N(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X ),
    .C(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X_sky130_fd_sc_hd__and3b_2_B_X ));
 sky130_fd_sc_hd__a31o_1 \prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1  (.A1(\prev2[10]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A3(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[12]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net77),
    .A2(net52),
    .B1(net60),
    .B2(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[12]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(\prev2[12]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[12] ));
 sky130_fd_sc_hd__nand2_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B  (.A(net76),
    .B(\prev2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A2(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__nand3_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .C(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__o21a_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1  (.A1(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(net82),
    .B1(\prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__o311a_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2  (.A1(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ),
    .A2(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .A3(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_A3 ),
    .B1(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_B1 ),
    .C1(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_C1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_X ));
 sky130_fd_sc_hd__nor2_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_A3_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev1[15] ),
    .B(\prev2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_A3 ));
 sky130_fd_sc_hd__nand3b_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_B1_sky130_fd_sc_hd__nand3b_2_Y  (.A_N(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_A3 ),
    .B(\prev2[14] ),
    .C(\prev1[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_B1 ));
 sky130_fd_sc_hd__nand2_1 \prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_C1_sky130_fd_sc_hd__nand2_2_Y  (.A(net86),
    .B(\prev2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o311a_2_A2_C1 ));
 sky130_fd_sc_hd__xnor2_1 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B  (.A(\prev1[12] ),
    .B(\prev2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__or2_4 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or2_2_A  (.A(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[12]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__or4_4 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A  (.A(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D ),
    .B(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .C(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ),
    .D(\prev2[13]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D_sky130_fd_sc_hd__xnor2_2_Y  (.A(\prev2[15] ),
    .B(\prev1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D ));
 sky130_fd_sc_hd__or3_4 \prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or3_2_C  (.A(\prev2[11]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ),
    .C(\prev2[10]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[13]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net75),
    .A2(net49),
    .B1(net57),
    .B2(\prev2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[13]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev2[13]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[13] ));
 sky130_fd_sc_hd__nand2_2 \prev2[13]_sky130_fd_sc_hd__nand2_2_B  (.A(net71),
    .B(\prev2[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__nand3_1 \prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\prev2[13]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev1[13]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .C(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__xnor2_4 \prev2[13]_sky130_fd_sc_hd__xnor2_2_B  (.A(\prev2[13] ),
    .B(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[13]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[14]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(\prev2[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[14] ));
 sky130_fd_sc_hd__a22o_1 \prev2[14]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\prev1[14] ),
    .A2(net49),
    .B1(net57),
    .B2(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[14]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_2 \prev2[14]_sky130_fd_sc_hd__xnor2_2_B  (.A(\prev1[14] ),
    .B(\prev2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_C ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[15]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev2[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[15] ));
 sky130_fd_sc_hd__a22o_1 \prev2[15]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(net84),
    .A2(net47),
    .B1(net55),
    .B2(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[15]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \prev2[16]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[16] ),
    .A2(net50),
    .B1(net59),
    .B2(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \prev2[16]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[16] ),
    .B(\prev2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[16]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \prev2[16]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A  (.A(\prev2[16]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_B1 ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[16]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(net133),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[16] ));
 sky130_fd_sc_hd__nor2_1 \prev2[16]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[16] ),
    .B(\prev2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\prev2[16]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\prev1[17] ),
    .A2(\prev2[17] ),
    .B1(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_B1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__inv_2 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A  (.A(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_4 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(net112),
    .B(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[18]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__o21bai_1 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A2  (.A1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A2(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1_N(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[20]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__o21a_1 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1  (.A1(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .A2(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_A2 ),
    .B1(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__o21ba_1 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1_sky130_fd_sc_hd__o21ba_2_X  (.A1(\prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1_N(\prev2[19]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_B1 ));
 sky130_fd_sc_hd__nor2_1 \prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A  (.A(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .B(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[17]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[17] ),
    .A2(net47),
    .B1(net55),
    .B2(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[17]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[17]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[17] ));
 sky130_fd_sc_hd__xor2_1 \prev2[17]_sky130_fd_sc_hd__xor2_2_B  (.A(\prev1[17] ),
    .B(\prev2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1  (.A1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1 ),
    .A2(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X ),
    .C1(\prev2[16]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[17]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__nand2_1 \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X_sky130_fd_sc_hd__and3b_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1 ));
 sky130_fd_sc_hd__nand2_1 \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[16]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21oi_4 \prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\prev2[11]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a211o_2_C1_X_sky130_fd_sc_hd__and3b_2_B_X ),
    .B1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[18]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net189),
    .A2(net47),
    .B1(net55),
    .B2(net146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[18]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[18]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[18] ));
 sky130_fd_sc_hd__nand2_1 \prev2[18]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[18] ),
    .B(\prev2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[18]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[18] ),
    .B(\prev2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[18]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or3_1 \prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\prev2[18]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev2[19]_sky130_fd_sc_hd__and2_2_B_X ),
    .C(\prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_A2 ));
 sky130_fd_sc_hd__a22o_1 \prev2[19]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[19] ),
    .A2(net46),
    .B1(net54),
    .B2(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \prev2[19]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[19] ),
    .B(\prev2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[19]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[19]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(net125),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[19] ));
 sky130_fd_sc_hd__nor2_1 \prev2[19]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[19] ),
    .B(\prev2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[19]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[1]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net103),
    .A2(net52),
    .B1(net60),
    .B2(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[1]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(net144),
    .RESET_B(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[1] ));
 sky130_fd_sc_hd__nand2_2 \prev2[1]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[1] ),
    .B(\prev2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[1]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_4 \prev2[1]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[1] ),
    .B(\prev2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21boi_2 \prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2  (.A1(\prev2[0]_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1_N(\prev2[1]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__a21o_1 \prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(\prev2[1]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\prev2[0]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[1]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__and3_1 \prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C  (.A(\prev2[0]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[1]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[20]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[20] ),
    .A2(net47),
    .B1(net55),
    .B2(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[20]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev2[20]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[20] ));
 sky130_fd_sc_hd__nand2_1 \prev2[20]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[20] ),
    .B(\prev2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[20]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[20] ),
    .B(\prev2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or3_1 \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_A2 ),
    .B(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2  (.A1(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A2(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[21]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[21] ),
    .A2(net46),
    .B1(net54),
    .B2(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[21]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(net130),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[21] ));
 sky130_fd_sc_hd__nand2_1 \prev2[21]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[21] ),
    .B(\prev2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[21] ),
    .B(\prev2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\prev2[20]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__a21oi_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\prev2[21]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__or4_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B  (.A(\prev2[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .C(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_C ),
    .D(\prev2[17]_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_C_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[21]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__or4_2_B_C ));
 sky130_fd_sc_hd__a22o_1 \prev2[22]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net192),
    .A2(net46),
    .B1(net54),
    .B2(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[22]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_0__leaf_clk),
    .D(\prev2[22]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[22] ));
 sky130_fd_sc_hd__nand2_1 \prev2[22]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[22] ),
    .B(\prev2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[22]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[22] ),
    .B(\prev2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[22]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or3_1 \prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev2[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .C(\prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[22]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[23]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[23] ),
    .A2(net46),
    .B1(net54),
    .B2(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \prev2[23]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[23] ),
    .B(\prev2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[23]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[23]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(net127),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[23] ));
 sky130_fd_sc_hd__nor2_1 \prev2[23]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[23] ),
    .B(\prev2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[23]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[24]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(\prev2[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[24] ));
 sky130_fd_sc_hd__a22o_1 \prev2[24]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\prev1[24] ),
    .A2(net46),
    .B1(net54),
    .B2(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[24]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \prev2[25]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[25] ),
    .A2(net48),
    .B1(net56),
    .B2(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[25]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_1__leaf_clk),
    .D(net142),
    .RESET_B(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[25] ));
 sky130_fd_sc_hd__nand2_1 \prev2[25]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[25] ),
    .B(\prev2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[25] ),
    .B(\prev2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A  (.A(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or4b_4 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4b_2_C  (.A(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .C(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .D_N(\prev2[20]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A ));
 sky130_fd_sc_hd__nand2b_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N ),
    .B(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A  (.A(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N ),
    .B(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__or2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__or2_2_X  (.A(\prev1[24] ),
    .B(\prev2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev1[24] ),
    .B(\prev2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_A_N ));
 sky130_fd_sc_hd__a211o_1 \prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2  (.A1(\prev2[25]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[25]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .C1(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_B1 ));
 sky130_fd_sc_hd__a22o_1 \prev2[26]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[26] ),
    .A2(net48),
    .B1(net56),
    .B2(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[26]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_4__leaf_clk),
    .D(net154),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[26] ));
 sky130_fd_sc_hd__nand2_1 \prev2[26]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[26] ),
    .B(\prev2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[26]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[26] ),
    .B(\prev2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[26]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[27]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[27] ),
    .A2(net49),
    .B1(net57),
    .B2(net160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[27]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev2[27]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[27] ));
 sky130_fd_sc_hd__nand2_1 \prev2[27]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[27] ),
    .B(\prev2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__inv_2 \prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__inv_2_A  (.A(\prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[27]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[27] ),
    .B(\prev2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211a_1 \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2  (.A1(\prev2[26]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_B1 ),
    .C1(\prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ));
 sky130_fd_sc_hd__a21oi_4 \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A ),
    .A2(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ),
    .B1(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__or3_2_X_A ));
 sky130_fd_sc_hd__nand2_4 \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__nand2_2_B  (.A(net85),
    .B(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ));
 sky130_fd_sc_hd__or2_1 \prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B  (.A(\prev2[27]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[28]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[28] ),
    .A2(net48),
    .B1(net56),
    .B2(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \prev2[28]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[28] ),
    .B(\prev2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1  (.A1(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ),
    .A2(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .C1(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[29]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__and2_1 \prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A  (.A(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[28]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(net148),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[28] ));
 sky130_fd_sc_hd__nor2_1 \prev2[28]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[28] ),
    .B(\prev2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[29]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net191),
    .A2(net48),
    .B1(net57),
    .B2(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \prev2[29]_sky130_fd_sc_hd__and2_2_B  (.A(\prev1[29] ),
    .B(\prev2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \prev2[29]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__or2_2_A  (.A(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\prev2[28]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__and2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[29]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev2[29]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[29] ));
 sky130_fd_sc_hd__nor2_1 \prev2[29]_sky130_fd_sc_hd__nor2_2_B  (.A(\prev1[29] ),
    .B(\prev2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\prev2[29]_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[28]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[29]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[2]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[2] ),
    .A2(net52),
    .B1(net61),
    .B2(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[2]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_6__leaf_clk),
    .D(net135),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[2] ));
 sky130_fd_sc_hd__nand2_1 \prev2[2]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[2] ),
    .B(\prev2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[2]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[2] ),
    .B(\prev2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[30]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[30] ),
    .A2(net48),
    .B1(net56),
    .B2(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[30]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(net138),
    .RESET_B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[30] ));
 sky130_fd_sc_hd__nand2_1 \prev2[30]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[30] ),
    .B(\prev2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[30]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[30]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[30] ),
    .B(\prev2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[30]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \prev2[30]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B  (.A(\prev2[30]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[30]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[30]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[31]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[31] ),
    .A2(net49),
    .B1(net57),
    .B2(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[31]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\prev2[31]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[31] ));
 sky130_fd_sc_hd__xnor2_1 \prev2[31]_sky130_fd_sc_hd__xnor2_2_B  (.A(\prev1[31] ),
    .B(\prev2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a21oi_2 \prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\prev2[30]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A1_N ));
 sky130_fd_sc_hd__a31o_1 \prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3  (.A1(\prev2[30]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev1[30]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .A3(\prev2[31]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B1(\iters[6]_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__nor2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[31]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a22o_1 \prev2[3]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net172),
    .A2(net50),
    .B1(net58),
    .B2(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[3]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev2[3]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[3] ));
 sky130_fd_sc_hd__nand2_1 \prev2[3]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[3] ),
    .B(\prev2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__o31a_1 \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1  (.A1(\prev2[1]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .A2(\prev2[2]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A3(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X ));
 sky130_fd_sc_hd__a211o_1 \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ),
    .A2(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B1(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B  (.A(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ),
    .B(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[4]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__or2_1 \prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__or2_2_X  (.A(\prev2[2]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__or2_1 \prev2[3]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[3] ),
    .B(\prev2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[3]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[4]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net193),
    .A2(net51),
    .B1(net58),
    .B2(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[4]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[4]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[4] ));
 sky130_fd_sc_hd__nand2_1 \prev2[4]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[4] ),
    .B(\prev2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[4]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[4] ),
    .B(\prev2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[4]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \prev2[5]_sky130_fd_sc_hd__a22o_2_B2  (.A1(net179),
    .A2(net51),
    .B1(net58),
    .B2(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[5]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[5]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[5] ));
 sky130_fd_sc_hd__nand2_2 \prev2[5]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[5] ),
    .B(\prev2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[5] ),
    .B(\prev2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_2 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or3_4 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__nand2b_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\prev2[4]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__a211o_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2  (.A1(\prev2[5]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ),
    .C1(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__o211a_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1  (.A1(\prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ),
    .B1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X ),
    .C1(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__nor2_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_A2_sky130_fd_sc_hd__nor2_2_Y  (.A(\prev1[7] ),
    .B(\prev2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ));
 sky130_fd_sc_hd__nand2_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1 ),
    .B(\prev2[7]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_A_C ));
 sky130_fd_sc_hd__nand2_1 \prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1_sky130_fd_sc_hd__nand2_2_Y  (.A(\prev1[7] ),
    .B(\prev2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[5]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a211o_2_A2_X_sky130_fd_sc_hd__o211a_2_B1_C1 ));
 sky130_fd_sc_hd__a22o_1 \prev2[6]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[6] ),
    .A2(net51),
    .B1(net58),
    .B2(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[6]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[6]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[6] ));
 sky130_fd_sc_hd__nand2_4 \prev2[6]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[6] ),
    .B(\prev2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_4 \prev2[6]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[6] ),
    .B(\prev2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_2 \prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A  (.A(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\prev2[6]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[6]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[7]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_2__leaf_clk),
    .D(\prev2[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[7] ));
 sky130_fd_sc_hd__a22o_1 \prev2[7]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\prev1[7] ),
    .A2(net50),
    .B1(net59),
    .B2(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[7]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \prev2[7]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[7] ),
    .B(\prev2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[7]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \prev2[8]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[8] ),
    .A2(net50),
    .B1(net59),
    .B2(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[8]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev2[8]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[8] ));
 sky130_fd_sc_hd__nand2_1 \prev2[8]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[8] ),
    .B(\prev2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[8]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[8] ),
    .B(\prev2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A  (.A(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a211o_4 \prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a211o_2_B1  (.A1(\prev2[3]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .A2(\prev1[8]_sky130_fd_sc_hd__dfrtp_2_Q_D_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X_B ),
    .B1(\prev2[8]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .C1(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or3_2_C_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__a211o_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__a22o_1 \prev2[9]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\prev1[9] ),
    .A2(net50),
    .B1(net59),
    .B2(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__dfrtp_1 \prev2[9]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_3__leaf_clk),
    .D(\prev2[9]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\prev2[9] ));
 sky130_fd_sc_hd__nand2_1 \prev2[9]_sky130_fd_sc_hd__nand2_2_B  (.A(\prev1[9] ),
    .B(\prev2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\prev2[8]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__nor2_2 \prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nor2_2_A  (.A(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .B(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or3_2_C_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \prev2[9]_sky130_fd_sc_hd__or2_2_B  (.A(\prev1[9] ),
    .B(\prev2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\prev2[9]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\prev2[9]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfstp_1 rdy_in_sky130_fd_sc_hd__dfstp_2_Q (.CLK(clknet_3_5__leaf_clk),
    .D(rdy_in_sky130_fd_sc_hd__dfstp_2_Q_D),
    .SET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net44));
 sky130_fd_sc_hd__a21bo_1 rdy_out_sky130_fd_sc_hd__a21bo_2_A2 (.A1(net159),
    .A2(net9),
    .B1_N(vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(rdy_in_sky130_fd_sc_hd__dfstp_2_Q_D));
 sky130_fd_sc_hd__o21ai_1 rdy_out_sky130_fd_sc_hd__o21ai_2_A2 (.A1(vld_out_sky130_fd_sc_hd__inv_2_A_Y),
    .A2(net9),
    .B1(rdy_out_sky130_fd_sc_hd__o21ai_2_A2_B1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(vld_out_sky130_fd_sc_hd__dfrtp_2_Q_D));
 sky130_fd_sc_hd__dfrtp_1 \state[2]_sky130_fd_sc_hd__dfrtp_2_Q  (.CLK(clknet_3_5__leaf_clk),
    .D(\state[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .RESET_B(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\state[2] ));
 sky130_fd_sc_hd__inv_2 \state[2]_sky130_fd_sc_hd__inv_2_A  (.A(\state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\state[2]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__or3_4 \state[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\state[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A1 ),
    .C(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(rdy_out_sky130_fd_sc_hd__o21ai_2_A2_B1));
 sky130_fd_sc_hd__o211ai_1 \state[2]_sky130_fd_sc_hd__o211ai_2_A1  (.A1(\state[2] ),
    .A2(net44),
    .B1(rdy_out_sky130_fd_sc_hd__o21ai_2_A2_B1),
    .C1(vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\state[2]_sky130_fd_sc_hd__o211ai_2_A1_Y ));
 sky130_fd_sc_hd__o21a_1 \state[2]_sky130_fd_sc_hd__o21a_2_B1  (.A1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A1 ),
    .A2(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A2 ),
    .B1(\state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and2_2_B  (.A(vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y),
    .B(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and3_2 \state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C  (.A(net64),
    .B(vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y),
    .C(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[0] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net121),
    .A1(net1),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[0]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[0] ),
    .B(\iters[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[1] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net116),
    .A1(net2),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[1]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[1] ),
    .B(\iters[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[2] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net117),
    .A1(net3),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[2]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[2] ),
    .B(\iters[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__or4_4 \target_iters[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A  (.A(\target_iters[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\target_iters[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .C(\target_iters[4]_sky130_fd_sc_hd__xor2_2_A_X ),
    .D(\target_iters[6]_sky130_fd_sc_hd__xor2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[3] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net115),
    .A1(net4),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[3]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[3] ),
    .B(\iters[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[3]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[4] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net119),
    .A1(net5),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[4]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[4] ),
    .B(\iters[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[4]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[5] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net114),
    .A1(net6),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[5]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[5] ),
    .B(\iters[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[6] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net122),
    .A1(net7),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[6]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[6] ),
    .B(\iters[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \target_iters[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_3_7__leaf_clk),
    .D(\target_iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\target_iters[7] ));
 sky130_fd_sc_hd__mux2_1 \target_iters[7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net118),
    .A1(net8),
    .S(vld_in_sky130_fd_sc_hd__and3_2_B_X),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \target_iters[7]_sky130_fd_sc_hd__xor2_2_A  (.A(\target_iters[7] ),
    .B(\iters[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\target_iters[7]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__or4_4 \target_iters[7]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A  (.A(\target_iters[7]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\target_iters[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .C(\target_iters[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .D(\target_iters[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__o21a_2_B1_A1 ));
 sky130_fd_sc_hd__a21o_1 vld_in_sky130_fd_sc_hd__a21o_2_A2 (.A1(net44),
    .A2(net11),
    .B1(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\state[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ));
 sky130_fd_sc_hd__and3_2 vld_in_sky130_fd_sc_hd__and3_2_B (.A(net44),
    .B(net11),
    .C(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(vld_in_sky130_fd_sc_hd__and3_2_B_X));
 sky130_fd_sc_hd__nand2b_1 vld_in_sky130_fd_sc_hd__nand2b_2_A_N (.A_N(net11),
    .B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(vld_in_sky130_fd_sc_hd__nand2b_2_A_N_Y));
 sky130_fd_sc_hd__dfrtp_1 vld_out_sky130_fd_sc_hd__dfrtp_2_Q (.CLK(clknet_3_5__leaf_clk),
    .D(vld_out_sky130_fd_sc_hd__dfrtp_2_Q_D),
    .RESET_B(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net45));
 sky130_fd_sc_hd__inv_2 vld_out_sky130_fd_sc_hd__inv_2_A (.A(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(vld_out_sky130_fd_sc_hd__inv_2_A_Y));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_74 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_76 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_77 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(fib_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(fib_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(fib_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(fib_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(fib_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(fib_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(fib_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(fib_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(rdy_out),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(vld_in),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[0]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[10]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[11]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[12]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[13]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[14]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[15]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[16]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[17]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[18]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[19]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[1]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[20]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[21]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[22]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[23]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[24]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[25]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[26]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[27]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[28]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[29]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[2]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[30]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[31]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[3]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[4]));
 sky130_fd_sc_hd__buf_6 output39 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[5]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[6]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[7]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[8]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(fib_out[9]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(rdy_in));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(vld_out));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(\state[2]_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__and2_2_B_X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 fanout59 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_6 fanout61 (.A(\state[2]_sky130_fd_sc_hd__o211ai_2_A1_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_4 clkload0 (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_4 clkload1 (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload5 (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer4 (.A(\prev1[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(\prev1[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(\prev1[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(\prev1[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(\prev2[13]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer15 (.A(\prev2[27]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer27 (.A(\prev1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(\prev2[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(\prev2[17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\target_iters[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\target_iters[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\target_iters[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\target_iters[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\target_iters[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\target_iters[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\target_iters[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\target_iters[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\prev2[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\prev2[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\prev2[19]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\prev2[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\prev2[23]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\prev2[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\prev2[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\prev2[21]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\prev2[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\prev2[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\prev2[16]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\prev2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\prev2[2]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\prev2[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\prev2[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\prev2[30]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\prev2[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\prev2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\prev2[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\prev2[25]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\prev2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\prev2[1]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\prev2[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\prev2[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\prev2[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\prev2[28]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\prev2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\prev2[0]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\prev2[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\iters[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\prev2[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\prev2[26]_sky130_fd_sc_hd__dfrtp_2_Q_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\prev2[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\prev2[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\iters[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\prev2[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\prev2[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\iters[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\prev2[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\prev2[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\prev2[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\prev2[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\prev1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\prev1[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\prev1[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\prev1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\prev1[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\prev1[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\prev1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\prev1[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\prev1[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\prev1[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\prev1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\prev1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\prev1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\prev1[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\prev1[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\prev1[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\prev1[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\prev1[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\prev1[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\prev2[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\prev2[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\iters[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\prev1[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\prev1[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\prev1[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\prev1[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\prev1[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\prev1[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(\prev1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(\prev1[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(\prev2[12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__or4_2_A_D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(\prev1[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(\prev1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_96 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_172 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_191 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_1_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_105 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_117 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_2_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_50 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_28 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_7_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_49 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_8_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_9_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_123 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_11_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_101 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_173 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_62 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_86 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_131 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_55 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_19_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_19_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_7 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_116 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_20_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_130 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_134 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_25_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_25_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_52 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_26_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_27_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_187 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_199 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_27_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_194 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_31_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_31_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_32_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_7 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_19 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_31 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_43 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_122 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_134 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_146 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_196 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_34_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_34_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_35_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
