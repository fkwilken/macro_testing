VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rcAdder
  CLASS BLOCK ;
  FOREIGN rcAdder ;
  ORIGIN 0.000 0.000 ;
  SIZE 62.115 BY 72.835 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 80.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 76.930 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 77.090 76.930 80.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.830 -9.470 76.930 80.190 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -9.470 25.940 80.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 30.030 76.930 31.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 75.390 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 72.130 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 72.290 72.130 75.390 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.030 -4.670 72.130 75.390 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -9.470 22.640 80.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 26.730 76.930 28.330 ;
    END
  END VPWR
  PIN a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 68.835 45.450 72.835 ;
    END
  END a_i[0]
  PIN a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END a_i[10]
  PIN a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END a_i[11]
  PIN a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END a_i[12]
  PIN a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END a_i[13]
  PIN a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END a_i[14]
  PIN a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END a_i[15]
  PIN a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 68.835 39.010 72.835 ;
    END
  END a_i[1]
  PIN a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 68.835 32.570 72.835 ;
    END
  END a_i[2]
  PIN a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 64.640 62.115 65.240 ;
    END
  END a_i[3]
  PIN a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 6.840 62.115 7.440 ;
    END
  END a_i[4]
  PIN a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 10.240 62.115 10.840 ;
    END
  END a_i[5]
  PIN a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 17.040 62.115 17.640 ;
    END
  END a_i[6]
  PIN a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END a_i[7]
  PIN a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END a_i[8]
  PIN a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END a_i[9]
  PIN b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.950 68.835 42.230 72.835 ;
    END
  END b_i[0]
  PIN b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END b_i[10]
  PIN b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b_i[11]
  PIN b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b_i[12]
  PIN b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END b_i[13]
  PIN b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END b_i[14]
  PIN b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END b_i[15]
  PIN b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.510 68.835 35.790 72.835 ;
    END
  END b_i[1]
  PIN b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 51.040 62.115 51.640 ;
    END
  END b_i[2]
  PIN b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 40.840 62.115 41.440 ;
    END
  END b_i[3]
  PIN b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 27.240 62.115 27.840 ;
    END
  END b_i[4]
  PIN b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 30.640 62.115 31.240 ;
    END
  END b_i[5]
  PIN b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 20.440 62.115 21.040 ;
    END
  END b_i[6]
  PIN b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END b_i[7]
  PIN b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END b_i[8]
  PIN b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END b_i[9]
  PIN carry_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END carry_o
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 58.115 61.240 62.115 61.840 ;
    END
  END clk
  PIN sum_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 57.840 62.115 58.440 ;
    END
  END sum_o[0]
  PIN sum_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END sum_o[10]
  PIN sum_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END sum_o[11]
  PIN sum_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END sum_o[12]
  PIN sum_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END sum_o[13]
  PIN sum_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 68.835 26.130 72.835 ;
    END
  END sum_o[14]
  PIN sum_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 68.835 29.350 72.835 ;
    END
  END sum_o[15]
  PIN sum_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 54.440 62.115 55.040 ;
    END
  END sum_o[1]
  PIN sum_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 47.640 62.115 48.240 ;
    END
  END sum_o[2]
  PIN sum_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 44.240 62.115 44.840 ;
    END
  END sum_o[3]
  PIN sum_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 34.040 62.115 34.640 ;
    END
  END sum_o[4]
  PIN sum_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 37.440 62.115 38.040 ;
    END
  END sum_o[5]
  PIN sum_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 23.840 62.115 24.440 ;
    END
  END sum_o[6]
  PIN sum_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 58.115 13.640 62.115 14.240 ;
    END
  END sum_o[7]
  PIN sum_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END sum_o[8]
  PIN sum_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END sum_o[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 56.770 59.925 ;
      LAYER li1 ;
        RECT 5.520 10.795 56.580 59.925 ;
      LAYER met1 ;
        RECT 4.210 10.640 56.580 60.080 ;
      LAYER met2 ;
        RECT 4.230 68.555 25.570 68.835 ;
        RECT 26.410 68.555 28.790 68.835 ;
        RECT 29.630 68.555 32.010 68.835 ;
        RECT 32.850 68.555 35.230 68.835 ;
        RECT 36.070 68.555 38.450 68.835 ;
        RECT 39.290 68.555 41.670 68.835 ;
        RECT 42.510 68.555 44.890 68.835 ;
        RECT 45.730 68.555 56.030 68.835 ;
        RECT 4.230 4.280 56.030 68.555 ;
        RECT 4.230 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 56.030 4.280 ;
      LAYER met3 ;
        RECT 4.400 64.240 57.715 65.105 ;
        RECT 3.990 62.240 58.115 64.240 ;
        RECT 4.400 60.840 57.715 62.240 ;
        RECT 3.990 58.840 58.115 60.840 ;
        RECT 4.400 57.440 57.715 58.840 ;
        RECT 3.990 55.440 58.115 57.440 ;
        RECT 4.400 54.040 57.715 55.440 ;
        RECT 3.990 52.040 58.115 54.040 ;
        RECT 4.400 50.640 57.715 52.040 ;
        RECT 3.990 48.640 58.115 50.640 ;
        RECT 4.400 47.240 57.715 48.640 ;
        RECT 3.990 45.240 58.115 47.240 ;
        RECT 4.400 43.840 57.715 45.240 ;
        RECT 3.990 41.840 58.115 43.840 ;
        RECT 4.400 40.440 57.715 41.840 ;
        RECT 3.990 38.440 58.115 40.440 ;
        RECT 4.400 37.040 57.715 38.440 ;
        RECT 3.990 35.040 58.115 37.040 ;
        RECT 4.400 33.640 57.715 35.040 ;
        RECT 3.990 31.640 58.115 33.640 ;
        RECT 4.400 30.240 57.715 31.640 ;
        RECT 3.990 28.240 58.115 30.240 ;
        RECT 4.400 26.840 57.715 28.240 ;
        RECT 3.990 24.840 58.115 26.840 ;
        RECT 4.400 23.440 57.715 24.840 ;
        RECT 3.990 21.440 58.115 23.440 ;
        RECT 4.400 20.040 57.715 21.440 ;
        RECT 3.990 18.040 58.115 20.040 ;
        RECT 4.400 16.640 57.715 18.040 ;
        RECT 3.990 14.640 58.115 16.640 ;
        RECT 3.990 13.240 57.715 14.640 ;
        RECT 3.990 11.240 58.115 13.240 ;
        RECT 3.990 9.840 57.715 11.240 ;
        RECT 3.990 7.840 58.115 9.840 ;
        RECT 3.990 6.975 57.715 7.840 ;
  END
END rcAdder
END LIBRARY

