magic
tech sky130A
magscale 1 2
timestamp 1740702134
<< viali >>
rect 1501 11849 1535 11883
rect 2329 11849 2363 11883
rect 2881 11849 2915 11883
rect 5457 11849 5491 11883
rect 6101 11849 6135 11883
rect 6469 11849 6503 11883
rect 7113 11849 7147 11883
rect 7757 11849 7791 11883
rect 8401 11849 8435 11883
rect 9045 11849 9079 11883
rect 3065 11781 3099 11815
rect 1685 11713 1719 11747
rect 1777 11713 1811 11747
rect 1961 11713 1995 11747
rect 2237 11713 2271 11747
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 5273 11713 5307 11747
rect 5917 11713 5951 11747
rect 6561 11713 6595 11747
rect 7205 11713 7239 11747
rect 8033 11713 8067 11747
rect 8493 11713 8527 11747
rect 9321 11713 9355 11747
rect 9965 11713 9999 11747
rect 10241 11713 10275 11747
rect 10609 11713 10643 11747
rect 10701 11713 10735 11747
rect 1961 11577 1995 11611
rect 2605 11577 2639 11611
rect 7849 11577 7883 11611
rect 10425 11577 10459 11611
rect 2053 11509 2087 11543
rect 3249 11509 3283 11543
rect 6745 11509 6779 11543
rect 7389 11509 7423 11543
rect 8677 11509 8711 11543
rect 9137 11509 9171 11543
rect 10057 11509 10091 11543
rect 10885 11509 10919 11543
rect 2237 11305 2271 11339
rect 5641 11305 5675 11339
rect 8677 11305 8711 11339
rect 10977 11305 11011 11339
rect 1501 11169 1535 11203
rect 2973 11169 3007 11203
rect 7205 11169 7239 11203
rect 7481 11169 7515 11203
rect 7757 11169 7791 11203
rect 8309 11169 8343 11203
rect 1685 11101 1719 11135
rect 1869 11101 1903 11135
rect 1961 11101 1995 11135
rect 2237 11101 2271 11135
rect 2421 11101 2455 11135
rect 2513 11101 2547 11135
rect 2697 11101 2731 11135
rect 3065 11101 3099 11135
rect 4261 11101 4295 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 7941 11101 7975 11135
rect 8033 11101 8067 11135
rect 8401 11101 8435 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9597 11101 9631 11135
rect 2605 11033 2639 11067
rect 4506 11033 4540 11067
rect 9842 11033 9876 11067
rect 3433 10965 3467 10999
rect 7573 10965 7607 10999
rect 8953 10965 8987 10999
rect 2421 10761 2455 10795
rect 5181 10761 5215 10795
rect 7665 10761 7699 10795
rect 8309 10761 8343 10795
rect 9137 10761 9171 10795
rect 10885 10761 10919 10795
rect 1869 10693 1903 10727
rect 9772 10693 9806 10727
rect 1409 10625 1443 10659
rect 1593 10625 1627 10659
rect 1685 10625 1719 10659
rect 2053 10625 2087 10659
rect 2513 10625 2547 10659
rect 2605 10625 2639 10659
rect 3801 10625 3835 10659
rect 4057 10625 4091 10659
rect 7021 10625 7055 10659
rect 7205 10625 7239 10659
rect 7389 10625 7423 10659
rect 7481 10625 7515 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 8769 10625 8803 10659
rect 8953 10625 8987 10659
rect 1501 10557 1535 10591
rect 2145 10557 2179 10591
rect 9505 10557 9539 10591
rect 6837 10421 6871 10455
rect 1685 10217 1719 10251
rect 3157 10217 3191 10251
rect 1961 10149 1995 10183
rect 8217 10149 8251 10183
rect 2789 10081 2823 10115
rect 6745 10081 6779 10115
rect 7205 10081 7239 10115
rect 7757 10081 7791 10115
rect 1409 10013 1443 10047
rect 1869 10013 1903 10047
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 2881 10013 2915 10047
rect 7113 10013 7147 10047
rect 7849 10013 7883 10047
rect 8125 10013 8159 10047
rect 8317 10013 8351 10047
rect 10333 10013 10367 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 2513 9945 2547 9979
rect 7389 9945 7423 9979
rect 1593 9877 1627 9911
rect 7481 9877 7515 9911
rect 10425 9877 10459 9911
rect 10885 9877 10919 9911
rect 1593 9605 1627 9639
rect 6561 9605 6595 9639
rect 6469 9537 6503 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 9873 9469 9907 9503
rect 8217 9401 8251 9435
rect 1409 9333 1443 9367
rect 9413 9333 9447 9367
rect 8677 9129 8711 9163
rect 2605 8993 2639 9027
rect 9229 8993 9263 9027
rect 9597 8993 9631 9027
rect 1409 8925 1443 8959
rect 1777 8925 1811 8959
rect 2145 8925 2179 8959
rect 2237 8925 2271 8959
rect 2421 8925 2455 8959
rect 2513 8925 2547 8959
rect 2697 8925 2731 8959
rect 7297 8925 7331 8959
rect 7564 8925 7598 8959
rect 9137 8925 9171 8959
rect 1961 8857 1995 8891
rect 9842 8857 9876 8891
rect 1593 8789 1627 8823
rect 2237 8789 2271 8823
rect 9505 8789 9539 8823
rect 10977 8789 11011 8823
rect 1961 8585 1995 8619
rect 2605 8585 2639 8619
rect 2789 8585 2823 8619
rect 9597 8585 9631 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 10057 8517 10091 8551
rect 1685 8449 1719 8483
rect 2329 8449 2363 8483
rect 3902 8449 3936 8483
rect 4169 8449 4203 8483
rect 9229 8449 9263 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 2421 8381 2455 8415
rect 9137 8381 9171 8415
rect 9873 8381 9907 8415
rect 1501 8313 1535 8347
rect 8953 8313 8987 8347
rect 10609 8041 10643 8075
rect 2605 7973 2639 8007
rect 2329 7905 2363 7939
rect 1685 7837 1719 7871
rect 2237 7837 2271 7871
rect 10701 7837 10735 7871
rect 1501 7701 1535 7735
rect 10885 7701 10919 7735
rect 2881 7497 2915 7531
rect 6929 7497 6963 7531
rect 8401 7497 8435 7531
rect 8217 7429 8251 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 3994 7361 4028 7395
rect 4261 7361 4295 7395
rect 9137 7361 9171 7395
rect 9393 7361 9427 7395
rect 10977 7361 11011 7395
rect 10517 7225 10551 7259
rect 1593 7157 1627 7191
rect 10793 7157 10827 7191
rect 2605 6953 2639 6987
rect 10977 6953 11011 6987
rect 3249 6885 3283 6919
rect 2421 6817 2455 6851
rect 2789 6817 2823 6851
rect 9045 6817 9079 6851
rect 1685 6749 1719 6783
rect 1869 6749 1903 6783
rect 2329 6749 2363 6783
rect 2881 6749 2915 6783
rect 9137 6749 9171 6783
rect 9597 6749 9631 6783
rect 1501 6681 1535 6715
rect 9842 6681 9876 6715
rect 1961 6613 1995 6647
rect 9505 6613 9539 6647
rect 1593 6409 1627 6443
rect 1961 6409 1995 6443
rect 2329 6409 2363 6443
rect 8493 6409 8527 6443
rect 9321 6409 9355 6443
rect 1409 6273 1443 6307
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 2145 6273 2179 6307
rect 2329 6273 2363 6307
rect 8125 6273 8159 6307
rect 8769 6273 8803 6307
rect 8861 6273 8895 6307
rect 9321 6273 9355 6307
rect 9505 6273 9539 6307
rect 10701 6273 10735 6307
rect 10977 6273 11011 6307
rect 8033 6205 8067 6239
rect 9229 6205 9263 6239
rect 8585 6069 8619 6103
rect 10793 6069 10827 6103
rect 1685 5865 1719 5899
rect 8217 5865 8251 5899
rect 9689 5865 9723 5899
rect 10241 5865 10275 5899
rect 10793 5797 10827 5831
rect 9413 5729 9447 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 8401 5661 8435 5695
rect 9321 5661 9355 5695
rect 9873 5661 9907 5695
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 10701 5661 10735 5695
rect 10977 5661 11011 5695
rect 8585 5593 8619 5627
rect 8769 5593 8803 5627
rect 10057 5593 10091 5627
rect 1593 5525 1627 5559
rect 8953 5525 8987 5559
rect 9597 5525 9631 5559
rect 2697 5321 2731 5355
rect 3341 5321 3375 5355
rect 8677 5321 8711 5355
rect 1777 5253 1811 5287
rect 3770 5253 3804 5287
rect 6745 5253 6779 5287
rect 1593 5185 1627 5219
rect 1961 5185 1995 5219
rect 2421 5185 2455 5219
rect 2973 5185 3007 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 10977 5185 11011 5219
rect 2053 5117 2087 5151
rect 2513 5117 2547 5151
rect 2881 5117 2915 5151
rect 3525 5117 3559 5151
rect 8493 5117 8527 5151
rect 4905 4981 4939 5015
rect 10793 4981 10827 5015
rect 1593 4777 1627 4811
rect 1869 4777 1903 4811
rect 2329 4777 2363 4811
rect 10977 4777 11011 4811
rect 9597 4641 9631 4675
rect 1409 4573 1443 4607
rect 1777 4573 1811 4607
rect 1961 4573 1995 4607
rect 2237 4573 2271 4607
rect 2421 4573 2455 4607
rect 2053 4505 2087 4539
rect 6745 4505 6779 4539
rect 9864 4505 9898 4539
rect 2881 4233 2915 4267
rect 9229 4233 9263 4267
rect 9873 4233 9907 4267
rect 10793 4233 10827 4267
rect 10425 4165 10459 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 4261 4097 4295 4131
rect 8861 4097 8895 4131
rect 9505 4097 9539 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 10241 4097 10275 4131
rect 10609 4097 10643 4131
rect 10977 4097 11011 4131
rect 2237 4029 2271 4063
rect 2605 4029 2639 4063
rect 2697 4029 2731 4063
rect 4169 4029 4203 4063
rect 8769 4029 8803 4063
rect 9413 4029 9447 4063
rect 10057 4029 10091 4063
rect 1593 3893 1627 3927
rect 4537 3893 4571 3927
rect 8585 3893 8619 3927
rect 1593 3689 1627 3723
rect 3801 3689 3835 3723
rect 4629 3689 4663 3723
rect 10241 3689 10275 3723
rect 10701 3689 10735 3723
rect 2145 3621 2179 3655
rect 10793 3621 10827 3655
rect 2329 3553 2363 3587
rect 4997 3553 5031 3587
rect 6837 3553 6871 3587
rect 9045 3553 9079 3587
rect 1501 3485 1535 3519
rect 1685 3485 1719 3519
rect 1961 3485 1995 3519
rect 2421 3485 2455 3519
rect 2881 3485 2915 3519
rect 3065 3485 3099 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 6469 3485 6503 3519
rect 6653 3485 6687 3519
rect 9137 3485 9171 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 1777 3417 1811 3451
rect 2973 3417 3007 3451
rect 5264 3417 5298 3451
rect 7082 3417 7116 3451
rect 2789 3349 2823 3383
rect 4445 3349 4479 3383
rect 6377 3349 6411 3383
rect 6561 3349 6595 3383
rect 8217 3349 8251 3383
rect 9505 3349 9539 3383
rect 1593 3145 1627 3179
rect 2697 3145 2731 3179
rect 4905 3145 4939 3179
rect 6101 3145 6135 3179
rect 6929 3145 6963 3179
rect 8769 3145 8803 3179
rect 3402 3077 3436 3111
rect 4997 3077 5031 3111
rect 9842 3077 9876 3111
rect 1409 3009 1443 3043
rect 1685 3009 1719 3043
rect 2881 3009 2915 3043
rect 3065 3009 3099 3043
rect 3157 3009 3191 3043
rect 4721 3009 4755 3043
rect 4905 3009 4939 3043
rect 5181 3009 5215 3043
rect 5641 3009 5675 3043
rect 6561 3009 6595 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 8309 3009 8343 3043
rect 8493 3009 8527 3043
rect 8585 3009 8619 3043
rect 8769 3009 8803 3043
rect 9597 3009 9631 3043
rect 5365 2941 5399 2975
rect 5733 2941 5767 2975
rect 6469 2941 6503 2975
rect 7389 2941 7423 2975
rect 8033 2941 8067 2975
rect 8125 2941 8159 2975
rect 4537 2873 4571 2907
rect 5457 2805 5491 2839
rect 10977 2805 11011 2839
rect 3065 2601 3099 2635
rect 3433 2601 3467 2635
rect 4813 2601 4847 2635
rect 5917 2601 5951 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 9137 2601 9171 2635
rect 10149 2601 10183 2635
rect 10425 2601 10459 2635
rect 10793 2601 10827 2635
rect 3985 2533 4019 2567
rect 2973 2397 3007 2431
rect 3249 2397 3283 2431
rect 3341 2397 3375 2431
rect 3525 2397 3559 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 6101 2397 6135 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 8125 2397 8159 2431
rect 8493 2397 8527 2431
rect 9321 2397 9355 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 10977 2397 11011 2431
rect 9873 2329 9907 2363
rect 3893 2261 3927 2295
rect 4537 2261 4571 2295
rect 5457 2261 5491 2295
rect 5825 2261 5859 2295
rect 6745 2261 6779 2295
rect 7389 2261 7423 2295
rect 7757 2261 7791 2295
rect 8677 2261 8711 2295
rect 9045 2261 9079 2295
<< metal1 >>
rect 1104 11994 11316 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 11316 11994
rect 1104 11920 11316 11942
rect 1026 11840 1032 11892
rect 1084 11880 1090 11892
rect 1489 11883 1547 11889
rect 1489 11880 1501 11883
rect 1084 11852 1501 11880
rect 1084 11840 1090 11852
rect 1489 11849 1501 11852
rect 1535 11849 1547 11883
rect 1489 11843 1547 11849
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 2332 11812 2360 11843
rect 2866 11840 2872 11892
rect 2924 11840 2930 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5316 11852 5457 11880
rect 5316 11840 5322 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 6089 11883 6147 11889
rect 6089 11880 6101 11883
rect 5868 11852 6101 11880
rect 5868 11840 5874 11852
rect 6089 11849 6101 11852
rect 6135 11849 6147 11883
rect 6089 11843 6147 11849
rect 6454 11840 6460 11892
rect 6512 11840 6518 11892
rect 7098 11840 7104 11892
rect 7156 11840 7162 11892
rect 7742 11840 7748 11892
rect 7800 11840 7806 11892
rect 8386 11840 8392 11892
rect 8444 11840 8450 11892
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 3053 11815 3111 11821
rect 3053 11812 3065 11815
rect 1780 11784 2360 11812
rect 2516 11784 3065 11812
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 1780 11753 1808 11784
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1780 11676 1808 11707
rect 1544 11648 1808 11676
rect 1544 11636 1550 11648
rect 1854 11636 1860 11688
rect 1912 11676 1918 11688
rect 1964 11676 1992 11707
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2188 11716 2237 11744
rect 2188 11704 2194 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2516 11753 2544 11784
rect 3053 11781 3065 11784
rect 3099 11781 3111 11815
rect 3053 11775 3111 11781
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 2372 11716 2513 11744
rect 2372 11704 2378 11716
rect 2501 11713 2513 11716
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 2866 11744 2872 11756
rect 2823 11716 2872 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5684 11716 5917 11744
rect 5684 11704 5690 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 6472 11744 6500 11840
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6472 11716 6561 11744
rect 5905 11707 5963 11713
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 7116 11744 7144 11840
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 7116 11716 7205 11744
rect 6549 11707 6607 11713
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7760 11744 7788 11840
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7760 11716 8033 11744
rect 7193 11707 7251 11713
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 8404 11744 8432 11840
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8404 11716 8493 11744
rect 8021 11707 8079 11713
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 9048 11744 9076 11840
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9048 11716 9321 11744
rect 8481 11707 8539 11713
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10226 11744 10232 11756
rect 9999 11716 10232 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 10686 11704 10692 11756
rect 10744 11704 10750 11756
rect 1912 11648 2636 11676
rect 1912 11636 1918 11648
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11608 2007 11611
rect 2406 11608 2412 11620
rect 1995 11580 2412 11608
rect 1995 11577 2007 11580
rect 1949 11571 2007 11577
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 2608 11617 2636 11648
rect 2593 11611 2651 11617
rect 2593 11577 2605 11611
rect 2639 11577 2651 11611
rect 2593 11571 2651 11577
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 7248 11580 7849 11608
rect 7248 11568 7254 11580
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7837 11571 7895 11577
rect 10410 11568 10416 11620
rect 10468 11568 10474 11620
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2041 11543 2099 11549
rect 2041 11540 2053 11543
rect 1820 11512 2053 11540
rect 1820 11500 1826 11512
rect 2041 11509 2053 11512
rect 2087 11509 2099 11543
rect 2041 11503 2099 11509
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 3237 11543 3295 11549
rect 3237 11540 3249 11543
rect 2188 11512 3249 11540
rect 2188 11500 2194 11512
rect 3237 11509 3249 11512
rect 3283 11509 3295 11543
rect 3237 11503 3295 11509
rect 6733 11543 6791 11549
rect 6733 11509 6745 11543
rect 6779 11540 6791 11543
rect 7098 11540 7104 11552
rect 6779 11512 7104 11540
rect 6779 11509 6791 11512
rect 6733 11503 6791 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7374 11500 7380 11552
rect 7432 11500 7438 11552
rect 8662 11500 8668 11552
rect 8720 11500 8726 11552
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 9306 11540 9312 11552
rect 9171 11512 9312 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 10134 11540 10140 11552
rect 10091 11512 10140 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 11146 11540 11152 11552
rect 10919 11512 11152 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 1104 11450 11316 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 11316 11450
rect 1104 11376 11316 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2225 11339 2283 11345
rect 2225 11336 2237 11339
rect 1728 11308 2237 11336
rect 1728 11296 1734 11308
rect 2225 11305 2237 11308
rect 2271 11305 2283 11339
rect 2225 11299 2283 11305
rect 5626 11296 5632 11348
rect 5684 11296 5690 11348
rect 8665 11339 8723 11345
rect 8665 11305 8677 11339
rect 8711 11336 8723 11339
rect 9766 11336 9772 11348
rect 8711 11308 9772 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10652 11308 10977 11336
rect 10652 11296 10658 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 1854 11228 1860 11280
rect 1912 11228 1918 11280
rect 2240 11240 3004 11268
rect 1486 11160 1492 11212
rect 1544 11160 1550 11212
rect 1872 11200 1900 11228
rect 1688 11172 1900 11200
rect 1688 11141 1716 11172
rect 2240 11144 2268 11240
rect 2976 11209 3004 11240
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 9306 11268 9312 11280
rect 7892 11240 9312 11268
rect 7892 11228 7898 11240
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 2961 11203 3019 11209
rect 2424 11172 2728 11200
rect 2424 11144 2452 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1903 11104 1961 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 1964 11064 1992 11095
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 2700 11141 2728 11172
rect 2961 11169 2973 11203
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7515 11172 7757 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 7745 11169 7757 11172
rect 7791 11200 7803 11203
rect 7791 11172 8156 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 2516 11064 2544 11095
rect 1964 11036 2544 11064
rect 2593 11067 2651 11073
rect 2593 11033 2605 11067
rect 2639 11064 2651 11067
rect 3068 11064 3096 11095
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 7006 11132 7012 11144
rect 4304 11104 7012 11132
rect 4304 11092 4310 11104
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7374 11132 7380 11144
rect 7147 11104 7380 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 4494 11067 4552 11073
rect 4494 11064 4506 11067
rect 2639 11036 3096 11064
rect 3436 11036 4506 11064
rect 2639 11033 2651 11036
rect 2593 11027 2651 11033
rect 3436 11005 3464 11036
rect 4494 11033 4506 11036
rect 4540 11033 4552 11067
rect 7944 11064 7972 11095
rect 8018 11092 8024 11144
rect 8076 11092 8082 11144
rect 8128 11132 8156 11172
rect 8294 11160 8300 11212
rect 8352 11160 8358 11212
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 8128 11104 8401 11132
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8720 11104 9137 11132
rect 8720 11092 8726 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9585 11135 9643 11141
rect 9585 11132 9597 11135
rect 9548 11104 9597 11132
rect 9548 11092 9554 11104
rect 9585 11101 9597 11104
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 8680 11064 8708 11092
rect 7944 11036 8708 11064
rect 4494 11027 4552 11033
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9830 11067 9888 11073
rect 9830 11064 9842 11067
rect 9732 11036 9842 11064
rect 9732 11024 9738 11036
rect 9830 11033 9842 11036
rect 9876 11033 9888 11067
rect 9830 11027 9888 11033
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10965 3479 10999
rect 3421 10959 3479 10965
rect 7558 10956 7564 11008
rect 7616 10956 7622 11008
rect 8938 10956 8944 11008
rect 8996 10956 9002 11008
rect 1104 10906 11316 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 11316 10906
rect 1104 10832 11316 10854
rect 1762 10792 1768 10804
rect 1504 10764 1768 10792
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1504 10656 1532 10764
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 2280 10764 2421 10792
rect 2280 10752 2286 10764
rect 2409 10761 2421 10764
rect 2455 10761 2467 10795
rect 2409 10755 2467 10761
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 7190 10752 7196 10804
rect 7248 10752 7254 10804
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 8018 10792 8024 10804
rect 7699 10764 8024 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9125 10795 9183 10801
rect 8352 10764 8800 10792
rect 8352 10752 8358 10764
rect 1857 10727 1915 10733
rect 1857 10724 1869 10727
rect 1596 10696 1869 10724
rect 1596 10668 1624 10696
rect 1857 10693 1869 10696
rect 1903 10693 1915 10727
rect 4246 10724 4252 10736
rect 1857 10687 1915 10693
rect 3804 10696 4252 10724
rect 1443 10628 1532 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1578 10616 1584 10668
rect 1636 10616 1642 10668
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1762 10656 1768 10668
rect 1719 10628 1768 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2498 10656 2504 10668
rect 2087 10628 2504 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 2682 10656 2688 10668
rect 2639 10628 2688 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3804 10665 3832 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 7208 10724 7236 10752
rect 7208 10696 7512 10724
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4045 10659 4103 10665
rect 4045 10656 4057 10659
rect 3936 10628 4057 10656
rect 3936 10616 3942 10628
rect 4045 10625 4057 10628
rect 4091 10625 4103 10659
rect 4045 10619 4103 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10588 1547 10591
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1535 10560 2145 10588
rect 1535 10557 1547 10560
rect 1489 10551 1547 10557
rect 2133 10557 2145 10560
rect 2179 10588 2191 10591
rect 2406 10588 2412 10600
rect 2179 10560 2412 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 7024 10588 7052 10619
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 7484 10665 7512 10696
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 7892 10628 8217 10656
rect 7892 10616 7898 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8662 10656 8668 10668
rect 8435 10628 8668 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8772 10665 8800 10764
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9674 10792 9680 10804
rect 9171 10764 9680 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10744 10764 10885 10792
rect 10744 10752 10750 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 9766 10733 9772 10736
rect 9760 10724 9772 10733
rect 9727 10696 9772 10724
rect 9760 10687 9772 10696
rect 9766 10684 9772 10687
rect 9824 10684 9830 10736
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 8294 10588 8300 10600
rect 7024 10560 8300 10588
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 9490 10548 9496 10600
rect 9548 10548 9554 10600
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 8110 10520 8116 10532
rect 7248 10492 8116 10520
rect 7248 10480 7254 10492
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 6822 10412 6828 10464
rect 6880 10412 6886 10464
rect 1104 10362 11316 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 11316 10362
rect 1104 10288 11316 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 1673 10251 1731 10257
rect 1673 10248 1685 10251
rect 1636 10220 1685 10248
rect 1636 10208 1642 10220
rect 1673 10217 1685 10220
rect 1719 10217 1731 10251
rect 1673 10211 1731 10217
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3878 10248 3884 10260
rect 3191 10220 3884 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 1302 10140 1308 10192
rect 1360 10180 1366 10192
rect 1949 10183 2007 10189
rect 1949 10180 1961 10183
rect 1360 10152 1961 10180
rect 1360 10140 1366 10152
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 1578 10044 1584 10056
rect 1443 10016 1584 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1872 10053 1900 10152
rect 1949 10149 1961 10152
rect 1995 10149 2007 10183
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 1949 10143 2007 10149
rect 6748 10152 8217 10180
rect 2498 10072 2504 10124
rect 2556 10072 2562 10124
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2740 10084 2789 10112
rect 2740 10072 2746 10084
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6748 10121 6776 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8205 10143 8263 10149
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6512 10084 6745 10112
rect 6512 10072 6518 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 6880 10084 7205 10112
rect 6880 10072 6886 10084
rect 7193 10081 7205 10084
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7742 10072 7748 10124
rect 7800 10072 7806 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 2516 10044 2544 10072
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 2516 10016 2605 10044
rect 2593 10013 2605 10016
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7558 10044 7564 10056
rect 7147 10016 7564 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9976 2559 9979
rect 2884 9976 2912 10007
rect 7558 10004 7564 10016
rect 7616 10044 7622 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7616 10016 7849 10044
rect 7616 10004 7622 10016
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8294 10004 8300 10056
rect 8352 10053 8358 10056
rect 8352 10044 8363 10053
rect 10321 10047 10379 10053
rect 8352 10016 9260 10044
rect 8352 10007 8363 10016
rect 8352 10004 8358 10007
rect 2547 9948 2912 9976
rect 7377 9979 7435 9985
rect 2547 9945 2559 9948
rect 2501 9939 2559 9945
rect 7377 9945 7389 9979
rect 7423 9976 7435 9979
rect 9122 9976 9128 9988
rect 7423 9948 9128 9976
rect 7423 9945 7435 9948
rect 7377 9939 7435 9945
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1762 9908 1768 9920
rect 1627 9880 1768 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 7558 9908 7564 9920
rect 7515 9880 7564 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 9232 9908 9260 10016
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 10594 10044 10600 10056
rect 10367 10016 10600 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 9232 9880 10425 9908
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 11146 9908 11152 9920
rect 10919 9880 11152 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 1104 9818 11316 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 11316 9818
rect 1104 9744 11316 9766
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 6549 9639 6607 9645
rect 6549 9605 6561 9639
rect 6595 9636 6607 9639
rect 7742 9636 7748 9648
rect 6595 9608 7748 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 10134 9636 10140 9648
rect 9784 9608 10140 9636
rect 6454 9528 6460 9580
rect 6512 9528 6518 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6822 9568 6828 9580
rect 6687 9540 6828 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9784 9577 9812 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10042 9568 10048 9580
rect 9999 9540 10048 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 9508 9500 9536 9531
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 9582 9500 9588 9512
rect 9508 9472 9588 9500
rect 9582 9460 9588 9472
rect 9640 9500 9646 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9640 9472 9873 9500
rect 9640 9460 9646 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7064 9404 8217 9432
rect 7064 9392 7070 9404
rect 8205 9401 8217 9404
rect 8251 9432 8263 9435
rect 9490 9432 9496 9444
rect 8251 9404 9496 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 1397 9367 1455 9373
rect 1397 9364 1409 9367
rect 1360 9336 1409 9364
rect 1360 9324 1366 9336
rect 1397 9333 1409 9336
rect 1443 9333 1455 9367
rect 1397 9327 1455 9333
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9272 9336 9413 9364
rect 9272 9324 9278 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 1104 9274 11316 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 11316 9274
rect 1104 9200 11316 9222
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 10686 9160 10692 9172
rect 8711 9132 10692 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 1762 9052 1768 9104
rect 1820 9092 1826 9104
rect 1820 9064 2728 9092
rect 1820 9052 1826 9064
rect 2593 9027 2651 9033
rect 2593 9024 2605 9027
rect 2424 8996 2605 9024
rect 2424 8968 2452 8996
rect 2593 8993 2605 8996
rect 2639 8993 2651 9027
rect 2593 8987 2651 8993
rect 1302 8916 1308 8968
rect 1360 8956 1366 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 1360 8928 1409 8956
rect 1360 8916 1366 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2179 8928 2237 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2225 8925 2237 8928
rect 2271 8956 2283 8959
rect 2314 8956 2320 8968
rect 2271 8928 2320 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 2406 8916 2412 8968
rect 2464 8916 2470 8968
rect 2700 8965 2728 9064
rect 9214 8984 9220 9036
rect 9272 8984 9278 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9548 8996 9597 9024
rect 9548 8984 9554 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9585 8987 9643 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 1949 8891 2007 8897
rect 1949 8857 1961 8891
rect 1995 8888 2007 8891
rect 2516 8888 2544 8919
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 7006 8956 7012 8968
rect 4212 8928 7012 8956
rect 4212 8916 4218 8928
rect 7006 8916 7012 8928
rect 7064 8956 7070 8968
rect 7558 8965 7564 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 7064 8928 7297 8956
rect 7064 8916 7070 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7552 8956 7564 8965
rect 7519 8928 7564 8956
rect 7285 8919 7343 8925
rect 7552 8919 7564 8928
rect 7558 8916 7564 8919
rect 7616 8916 7622 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9830 8891 9888 8897
rect 9830 8888 9842 8891
rect 1995 8860 2544 8888
rect 9508 8860 9842 8888
rect 1995 8857 2007 8860
rect 1949 8851 2007 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1964 8820 1992 8851
rect 1627 8792 1992 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 2222 8780 2228 8832
rect 2280 8780 2286 8832
rect 9508 8829 9536 8860
rect 9830 8857 9842 8860
rect 9876 8857 9888 8891
rect 9830 8851 9888 8857
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8789 9551 8823
rect 9493 8783 9551 8789
rect 10962 8780 10968 8832
rect 11020 8780 11026 8832
rect 1104 8730 11316 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 11316 8730
rect 1104 8656 11316 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2406 8616 2412 8628
rect 1995 8588 2412 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2593 8619 2651 8625
rect 2593 8585 2605 8619
rect 2639 8616 2651 8619
rect 2682 8616 2688 8628
rect 2639 8588 2688 8616
rect 2639 8585 2651 8588
rect 2593 8579 2651 8585
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8585 2835 8619
rect 2777 8579 2835 8585
rect 2792 8548 2820 8579
rect 9582 8576 9588 8628
rect 9640 8576 9646 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 1688 8520 2820 8548
rect 1688 8489 1716 8520
rect 9122 8508 9128 8560
rect 9180 8548 9186 8560
rect 9180 8520 9260 8548
rect 9180 8508 9186 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3890 8483 3948 8489
rect 3890 8480 3902 8483
rect 2832 8452 3902 8480
rect 2832 8440 2838 8452
rect 3890 8449 3902 8452
rect 3936 8449 3948 8483
rect 3890 8443 3948 8449
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 9232 8489 9260 8520
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 10428 8548 10456 8579
rect 10778 8576 10784 8628
rect 10836 8576 10842 8628
rect 10100 8520 10456 8548
rect 10100 8508 10106 8520
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 10192 8452 10241 8480
rect 10192 8440 10198 8452
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8381 2467 8415
rect 2409 8375 2467 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9306 8412 9312 8424
rect 9171 8384 9312 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2424 8344 2452 8375
rect 9306 8372 9312 8384
rect 9364 8412 9370 8424
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 9364 8384 9873 8412
rect 9364 8372 9370 8384
rect 9861 8381 9873 8384
rect 9907 8381 9919 8415
rect 9861 8375 9919 8381
rect 2372 8316 2452 8344
rect 8941 8347 8999 8353
rect 2372 8304 2378 8316
rect 8941 8313 8953 8347
rect 8987 8344 8999 8347
rect 9030 8344 9036 8356
rect 8987 8316 9036 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 1104 8186 11316 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 11316 8186
rect 1104 8112 11316 8134
rect 10594 8032 10600 8084
rect 10652 8032 10658 8084
rect 2593 8007 2651 8013
rect 2593 7973 2605 8007
rect 2639 8004 2651 8007
rect 2774 8004 2780 8016
rect 2639 7976 2780 8004
rect 2639 7973 2651 7976
rect 2593 7967 2651 7973
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 2314 7896 2320 7948
rect 2372 7896 2378 7948
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10560 7840 10701 7868
rect 10560 7828 10566 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 10870 7692 10876 7744
rect 10928 7692 10934 7744
rect 1104 7642 11316 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 11316 7642
rect 1104 7568 11316 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 1728 7500 2881 7528
rect 1728 7488 1734 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 8220 7500 8401 7528
rect 8220 7469 8248 7500
rect 8389 7497 8401 7500
rect 8435 7528 8447 7531
rect 11054 7528 11060 7540
rect 8435 7500 11060 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7429 8263 7463
rect 9490 7460 9496 7472
rect 8205 7423 8263 7429
rect 9140 7432 9496 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1360 7364 1409 7392
rect 1360 7352 1366 7364
rect 1397 7361 1409 7364
rect 1443 7392 1455 7395
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1443 7364 1685 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3982 7395 4040 7401
rect 3982 7392 3994 7395
rect 3292 7364 3994 7392
rect 3292 7352 3298 7364
rect 3982 7361 3994 7364
rect 4028 7361 4040 7395
rect 3982 7355 4040 7361
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 9140 7401 9168 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4212 7364 4261 7392
rect 4212 7352 4218 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9381 7395 9439 7401
rect 9381 7392 9393 7395
rect 9272 7364 9393 7392
rect 9272 7352 9278 7364
rect 9381 7361 9393 7364
rect 9427 7361 9439 7395
rect 9381 7355 9439 7361
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 10502 7216 10508 7268
rect 10560 7216 10566 7268
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11054 7188 11060 7200
rect 10827 7160 11060 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 1104 7098 11316 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 11316 7098
rect 1104 7024 11316 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2593 6987 2651 6993
rect 2593 6984 2605 6987
rect 2372 6956 2605 6984
rect 2372 6944 2378 6956
rect 2593 6953 2605 6956
rect 2639 6953 2651 6987
rect 2593 6947 2651 6953
rect 10962 6944 10968 6996
rect 11020 6944 11026 6996
rect 3234 6876 3240 6928
rect 3292 6876 3298 6928
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2682 6848 2688 6860
rect 2455 6820 2688 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2682 6808 2688 6820
rect 2740 6848 2746 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2740 6820 2789 6848
rect 2740 6808 2746 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9030 6848 9036 6860
rect 8812 6820 9036 6848
rect 8812 6808 8818 6820
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 2314 6780 2320 6792
rect 1903 6752 2320 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 2866 6740 2872 6792
rect 2924 6740 2930 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9306 6780 9312 6792
rect 9171 6752 9312 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 1489 6715 1547 6721
rect 1489 6681 1501 6715
rect 1535 6712 1547 6715
rect 1578 6712 1584 6724
rect 1535 6684 1584 6712
rect 1535 6681 1547 6684
rect 1489 6675 1547 6681
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 9830 6715 9888 6721
rect 9830 6712 9842 6715
rect 9508 6684 9842 6712
rect 1946 6604 1952 6656
rect 2004 6604 2010 6656
rect 9508 6653 9536 6684
rect 9830 6681 9842 6684
rect 9876 6681 9888 6715
rect 9830 6675 9888 6681
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6613 9551 6647
rect 9493 6607 9551 6613
rect 1104 6554 11316 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 11316 6554
rect 1104 6480 11316 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 1946 6400 1952 6452
rect 2004 6400 2010 6452
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2866 6440 2872 6452
rect 2363 6412 2872 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 9214 6440 9220 6452
rect 8527 6412 9220 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 1360 6276 1409 6304
rect 1360 6264 1366 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1596 6304 1624 6400
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 1964 6372 1992 6400
rect 1728 6344 1900 6372
rect 1964 6344 2176 6372
rect 1728 6332 1734 6344
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1596 6276 1777 6304
rect 1397 6267 1455 6273
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1872 6304 1900 6344
rect 2148 6313 2176 6344
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1872 6276 1961 6304
rect 1765 6267 1823 6273
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8202 6304 8208 6316
rect 8159 6276 8208 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 9306 6304 9312 6316
rect 8895 6276 9312 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 10226 6304 10232 6316
rect 9539 6276 10232 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 9217 6239 9275 6245
rect 8067 6208 8616 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 8588 6112 8616 6208
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 9508 6236 9536 6267
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10962 6304 10968 6316
rect 10735 6276 10968 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 9263 6208 9536 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 8720 6072 10793 6100
rect 8720 6060 8726 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 1104 6010 11316 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 11316 6010
rect 1104 5936 11316 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 1673 5899 1731 5905
rect 1673 5896 1685 5899
rect 1360 5868 1685 5896
rect 1360 5856 1366 5868
rect 1673 5865 1685 5868
rect 1719 5865 1731 5899
rect 1673 5859 1731 5865
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 9364 5868 9689 5896
rect 9364 5856 9370 5868
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 10226 5856 10232 5908
rect 10284 5856 10290 5908
rect 10781 5831 10839 5837
rect 10781 5797 10793 5831
rect 10827 5797 10839 5831
rect 10781 5791 10839 5797
rect 8128 5732 8432 5760
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 8128 5701 8156 5732
rect 8404 5701 8432 5732
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 8628 5732 9413 5760
rect 8628 5720 8634 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 10796 5760 10824 5791
rect 9401 5723 9459 5729
rect 10152 5732 10824 5760
rect 10152 5701 10180 5732
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1452 5664 1869 5692
rect 1452 5652 1458 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 8435 5664 9321 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9907 5664 10149 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10410 5692 10416 5704
rect 10367 5664 10416 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1762 5556 1768 5568
rect 1627 5528 1768 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 8312 5556 8340 5655
rect 8570 5584 8576 5636
rect 8628 5584 8634 5636
rect 8754 5584 8760 5636
rect 8812 5584 8818 5636
rect 10045 5627 10103 5633
rect 10045 5593 10057 5627
rect 10091 5624 10103 5627
rect 10336 5624 10364 5655
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10735 5664 10977 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 10965 5661 10977 5664
rect 11011 5692 11023 5695
rect 11146 5692 11152 5704
rect 11011 5664 11152 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 10091 5596 10364 5624
rect 10091 5593 10103 5596
rect 10045 5587 10103 5593
rect 8662 5556 8668 5568
rect 8312 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5556 8726 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8720 5528 8953 5556
rect 8720 5516 8726 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 8941 5519 8999 5525
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 9585 5559 9643 5565
rect 9585 5556 9597 5559
rect 9456 5528 9597 5556
rect 9456 5516 9462 5528
rect 9585 5525 9597 5528
rect 9631 5525 9643 5559
rect 9585 5519 9643 5525
rect 1104 5466 11316 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 11316 5466
rect 1104 5392 11316 5414
rect 2682 5312 2688 5364
rect 2740 5312 2746 5364
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5321 3387 5355
rect 3329 5315 3387 5321
rect 1762 5244 1768 5296
rect 1820 5244 1826 5296
rect 3344 5284 3372 5315
rect 8662 5312 8668 5364
rect 8720 5312 8726 5364
rect 3758 5287 3816 5293
rect 3758 5284 3770 5287
rect 3344 5256 3770 5284
rect 3758 5253 3770 5256
rect 3804 5253 3816 5287
rect 3758 5247 3816 5253
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 6914 5284 6920 5296
rect 6779 5256 6920 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2406 5216 2412 5228
rect 1995 5188 2412 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2958 5176 2964 5228
rect 3016 5176 3022 5228
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9674 5216 9680 5228
rect 8812 5188 9680 5216
rect 8812 5176 8818 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 1912 5120 2053 5148
rect 1912 5108 1918 5120
rect 2041 5117 2053 5120
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2866 5148 2872 5160
rect 2547 5120 2872 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3510 5108 3516 5160
rect 3568 5108 3574 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 6788 5120 8493 5148
rect 6788 5108 6794 5120
rect 8481 5117 8493 5120
rect 8527 5148 8539 5151
rect 9582 5148 9588 5160
rect 8527 5120 9588 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4856 4984 4905 5012
rect 4856 4972 4862 4984
rect 4893 4981 4905 4984
rect 4939 4981 4951 5015
rect 4893 4975 4951 4981
rect 10778 4972 10784 5024
rect 10836 4972 10842 5024
rect 1104 4922 11316 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 11316 4922
rect 1104 4848 11316 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 1854 4768 1860 4820
rect 1912 4768 1918 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2958 4808 2964 4820
rect 2363 4780 2964 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 10962 4768 10968 4820
rect 11020 4768 11026 4820
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 1360 4576 1409 4604
rect 1360 4564 1366 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1596 4604 1624 4768
rect 1872 4672 1900 4768
rect 1872 4644 2268 4672
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1596 4576 1777 4604
rect 1397 4567 1455 4573
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 1412 4536 1440 4567
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2240 4613 2268 4644
rect 9582 4632 9588 4684
rect 9640 4632 9646 4684
rect 1949 4607 2007 4613
rect 1949 4604 1961 4607
rect 1912 4576 1961 4604
rect 1912 4564 1918 4576
rect 1949 4573 1961 4576
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2406 4564 2412 4616
rect 2464 4564 2470 4616
rect 2041 4539 2099 4545
rect 2041 4536 2053 4539
rect 1412 4508 2053 4536
rect 2041 4505 2053 4508
rect 2087 4505 2099 4539
rect 2041 4499 2099 4505
rect 6730 4496 6736 4548
rect 6788 4496 6794 4548
rect 9858 4545 9864 4548
rect 9852 4499 9864 4545
rect 9858 4496 9864 4499
rect 9916 4496 9922 4548
rect 1104 4378 11316 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 11316 4378
rect 1104 4304 11316 4326
rect 2866 4224 2872 4276
rect 2924 4224 2930 4276
rect 9217 4267 9275 4273
rect 9217 4233 9229 4267
rect 9263 4264 9275 4267
rect 9263 4236 9812 4264
rect 9263 4233 9275 4236
rect 9217 4227 9275 4233
rect 9784 4196 9812 4236
rect 9858 4224 9864 4276
rect 9916 4224 9922 4276
rect 10134 4264 10140 4276
rect 9968 4236 10140 4264
rect 9968 4196 9996 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10428 4236 10793 4264
rect 9416 4168 9628 4196
rect 9784 4168 9996 4196
rect 10060 4168 10272 4196
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 1268 4100 1409 4128
rect 1268 4088 1274 4100
rect 1397 4097 1409 4100
rect 1443 4128 1455 4131
rect 1673 4131 1731 4137
rect 1673 4128 1685 4131
rect 1443 4100 1685 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1673 4097 1685 4100
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4614 4128 4620 4140
rect 4295 4100 4620 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9416 4128 9444 4168
rect 8895 4100 9444 4128
rect 9493 4131 9551 4137
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9600 4128 9628 4168
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9600 4100 9965 4128
rect 9493 4091 9551 4097
rect 9953 4097 9965 4100
rect 9999 4128 10011 4131
rect 10060 4128 10088 4168
rect 9999 4100 10088 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 1636 4032 2237 4060
rect 1636 4020 1642 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2240 3992 2268 4023
rect 2590 4020 2596 4072
rect 2648 4020 2654 4072
rect 2682 4020 2688 4072
rect 2740 4020 2746 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 4120 4032 4169 4060
rect 4120 4020 4126 4032
rect 4157 4029 4169 4032
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 3050 3992 3056 4004
rect 2240 3964 3056 3992
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 8772 3992 8800 4023
rect 9398 4020 9404 4072
rect 9456 4020 9462 4072
rect 9508 4060 9536 4091
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 10244 4137 10272 4168
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 10428 4205 10456 4236
rect 10781 4233 10793 4236
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 10413 4199 10471 4205
rect 10413 4196 10425 4199
rect 10376 4168 10425 4196
rect 10376 4156 10382 4168
rect 10413 4165 10425 4168
rect 10459 4165 10471 4199
rect 10413 4159 10471 4165
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10778 4128 10784 4140
rect 10643 4100 10784 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10962 4088 10968 4140
rect 11020 4088 11026 4140
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9508 4032 10057 4060
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 9416 3992 9444 4020
rect 8772 3964 9444 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1670 3924 1676 3936
rect 1627 3896 1676 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 5258 3924 5264 3936
rect 4571 3896 5264 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 7616 3896 8585 3924
rect 7616 3884 7622 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 1104 3834 11316 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 11316 3834
rect 1104 3760 11316 3782
rect 1578 3680 1584 3732
rect 1636 3680 1642 3732
rect 2682 3720 2688 3732
rect 2056 3692 2688 3720
rect 2056 3584 2084 3692
rect 2682 3680 2688 3692
rect 2740 3720 2746 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 2740 3692 3801 3720
rect 2740 3680 2746 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 4614 3680 4620 3732
rect 4672 3680 4678 3732
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10192 3692 10241 3720
rect 10192 3680 10198 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10962 3720 10968 3732
rect 10735 3692 10968 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 2133 3655 2191 3661
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2590 3652 2596 3664
rect 2179 3624 2596 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 2590 3612 2596 3624
rect 2648 3652 2654 3664
rect 2648 3624 2912 3652
rect 2648 3612 2654 3624
rect 2317 3587 2375 3593
rect 2317 3584 2329 3587
rect 2056 3556 2329 3584
rect 2317 3553 2329 3556
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 1486 3476 1492 3528
rect 1544 3476 1550 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2884 3525 2912 3624
rect 10778 3612 10784 3664
rect 10836 3612 10842 3664
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3510 3584 3516 3596
rect 3200 3556 3516 3584
rect 3200 3544 3206 3556
rect 3510 3544 3516 3556
rect 3568 3584 3574 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 3568 3556 4997 3584
rect 3568 3544 3574 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 6730 3584 6736 3596
rect 4985 3547 5043 3553
rect 6380 3556 6736 3584
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1728 3488 1961 3516
rect 1728 3476 1734 3488
rect 1949 3485 1961 3488
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 1504 3448 1532 3476
rect 1765 3451 1823 3457
rect 1765 3448 1777 3451
rect 1504 3420 1777 3448
rect 1765 3417 1777 3420
rect 1811 3417 1823 3451
rect 2424 3448 2452 3479
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 2961 3451 3019 3457
rect 2961 3448 2973 3451
rect 2424 3420 2973 3448
rect 1765 3411 1823 3417
rect 2961 3417 2973 3420
rect 3007 3417 3019 3451
rect 3988 3448 4016 3479
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4120 3488 4537 3516
rect 4120 3476 4126 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4525 3479 4583 3485
rect 4632 3488 4721 3516
rect 4154 3448 4160 3460
rect 3988 3420 4160 3448
rect 2961 3411 3019 3417
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4632 3392 4660 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 5000 3516 5028 3547
rect 6380 3516 6408 3556
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6788 3556 6837 3584
rect 6788 3544 6794 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 6825 3547 6883 3553
rect 8404 3556 9045 3584
rect 5000 3488 6408 3516
rect 4709 3479 4767 3485
rect 6454 3476 6460 3528
rect 6512 3476 6518 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 5258 3457 5264 3460
rect 5252 3448 5264 3457
rect 5219 3420 5264 3448
rect 5252 3411 5264 3420
rect 5258 3408 5264 3411
rect 5316 3408 5322 3460
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6656 3448 6684 3479
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 8404 3516 8432 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 10796 3584 10824 3612
rect 9033 3547 9091 3553
rect 10152 3556 10824 3584
rect 7616 3488 8432 3516
rect 7616 3476 7622 3488
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10152 3525 10180 3556
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8812 3488 9137 3516
rect 8812 3476 8818 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10318 3476 10324 3528
rect 10376 3476 10382 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10962 3516 10968 3528
rect 10551 3488 10968 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 5776 3420 6684 3448
rect 5776 3408 5782 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7070 3451 7128 3457
rect 7070 3448 7082 3451
rect 6972 3420 7082 3448
rect 6972 3408 6978 3420
rect 7070 3417 7082 3420
rect 7116 3417 7128 3451
rect 7070 3411 7128 3417
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4614 3380 4620 3392
rect 4479 3352 4620 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 6362 3340 6368 3392
rect 6420 3340 6426 3392
rect 6546 3340 6552 3392
rect 6604 3340 6610 3392
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8478 3380 8484 3392
rect 8251 3352 8484 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 9490 3340 9496 3392
rect 9548 3340 9554 3392
rect 1104 3290 11316 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 11316 3290
rect 1104 3216 11316 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 4062 3176 4068 3188
rect 2731 3148 4068 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 4939 3148 6101 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 6089 3145 6101 3148
rect 6135 3176 6147 3179
rect 6454 3176 6460 3188
rect 6135 3148 6460 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 3390 3111 3448 3117
rect 3390 3108 3402 3111
rect 2832 3080 3402 3108
rect 2832 3068 2838 3080
rect 3390 3077 3402 3080
rect 3436 3077 3448 3111
rect 4985 3111 5043 3117
rect 4985 3108 4997 3111
rect 3390 3071 3448 3077
rect 4724 3080 4997 3108
rect 4724 3052 4752 3080
rect 4985 3077 4997 3080
rect 5031 3077 5043 3111
rect 4985 3071 5043 3077
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8076 3080 8616 3108
rect 8076 3068 8082 3080
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1360 3012 1409 3040
rect 1360 3000 1366 3012
rect 1397 3009 1409 3012
rect 1443 3040 1455 3043
rect 1673 3043 1731 3049
rect 1673 3040 1685 3043
rect 1443 3012 1685 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1673 3009 1685 3012
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3142 3000 3148 3052
rect 3200 3000 3206 3052
rect 4706 3000 4712 3052
rect 4764 3000 4770 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 4939 3012 5181 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5169 3009 5181 3012
rect 5215 3040 5227 3043
rect 5534 3040 5540 3052
rect 5215 3012 5540 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5675 3012 6500 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2972 5411 2975
rect 5718 2972 5724 2984
rect 5399 2944 5724 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 6472 2981 6500 3012
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7699 3012 8156 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2972 6515 2975
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6503 2944 7389 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 8018 2932 8024 2984
rect 8076 2932 8082 2984
rect 8128 2981 8156 3012
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8588 3049 8616 3080
rect 9490 3068 9496 3120
rect 9548 3108 9554 3120
rect 9830 3111 9888 3117
rect 9830 3108 9842 3111
rect 9548 3080 9842 3108
rect 9548 3068 9554 3080
rect 9830 3077 9842 3080
rect 9876 3077 9888 3111
rect 9830 3071 9888 3077
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8444 3012 8493 3040
rect 8444 3000 8450 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 8772 2972 8800 3003
rect 9582 3000 9588 3052
rect 9640 3000 9646 3052
rect 8159 2944 8800 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2904 4583 2907
rect 7190 2904 7196 2916
rect 4571 2876 7196 2904
rect 4571 2873 4583 2876
rect 4525 2867 4583 2873
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 5445 2839 5503 2845
rect 5445 2836 5457 2839
rect 4212 2808 5457 2836
rect 4212 2796 4218 2808
rect 5445 2805 5457 2808
rect 5491 2805 5503 2839
rect 5445 2799 5503 2805
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 1104 2746 11316 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 11316 2746
rect 1104 2672 11316 2694
rect 3050 2592 3056 2644
rect 3108 2592 3114 2644
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 4614 2632 4620 2644
rect 3467 2604 4620 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4764 2604 4813 2632
rect 4764 2592 4770 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 4801 2595 4859 2601
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5592 2604 5917 2632
rect 5592 2592 5598 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 5905 2595 5963 2601
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8018 2632 8024 2644
rect 7975 2604 8024 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8294 2592 8300 2644
rect 8352 2592 8358 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8444 2604 9137 2632
rect 8444 2592 8450 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 9732 2604 10149 2632
rect 9732 2592 9738 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11054 2632 11060 2644
rect 10827 2604 11060 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 3068 2496 3096 2592
rect 3973 2567 4031 2573
rect 3973 2564 3985 2567
rect 3528 2536 3985 2564
rect 3068 2468 3372 2496
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3234 2428 3240 2440
rect 3007 2400 3240 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3344 2437 3372 2468
rect 3528 2437 3556 2536
rect 3973 2533 3985 2536
rect 4019 2533 4031 2567
rect 8202 2564 8208 2576
rect 3973 2527 4031 2533
rect 7852 2536 8208 2564
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 3513 2391 3571 2397
rect 3896 2400 4169 2428
rect 2866 2320 2872 2372
rect 2924 2360 2930 2372
rect 3528 2360 3556 2391
rect 2924 2332 3556 2360
rect 2924 2320 2930 2332
rect 3896 2304 3924 2400
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4157 2391 4215 2397
rect 4540 2400 4629 2428
rect 4540 2304 4568 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4856 2400 5273 2428
rect 4856 2388 4862 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5261 2391 5319 2397
rect 5828 2400 6101 2428
rect 5828 2304 5856 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7852 2437 7880 2536
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 8312 2496 8340 2592
rect 8036 2468 8340 2496
rect 8036 2437 8064 2468
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8128 2360 8156 2391
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9048 2400 9321 2428
rect 7760 2332 8156 2360
rect 7760 2304 7788 2332
rect 9048 2304 9076 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10318 2428 10324 2440
rect 10091 2400 10324 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 10962 2388 10968 2440
rect 11020 2388 11026 2440
rect 9861 2363 9919 2369
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 10612 2360 10640 2388
rect 9907 2332 10640 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 3878 2252 3884 2304
rect 3936 2252 3942 2304
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5316 2264 5457 2292
rect 5316 2252 5322 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8444 2264 8677 2292
rect 8444 2252 8450 2264
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 9030 2252 9036 2304
rect 9088 2252 9094 2304
rect 1104 2202 11316 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 11316 2202
rect 1104 2128 11316 2150
<< via1 >>
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 1032 11840 1084 11892
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 5264 11840 5316 11892
rect 5816 11840 5868 11892
rect 6460 11883 6512 11892
rect 6460 11849 6469 11883
rect 6469 11849 6503 11883
rect 6503 11849 6512 11883
rect 6460 11840 6512 11849
rect 7104 11883 7156 11892
rect 7104 11849 7113 11883
rect 7113 11849 7147 11883
rect 7147 11849 7156 11883
rect 7104 11840 7156 11849
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 8392 11883 8444 11892
rect 8392 11849 8401 11883
rect 8401 11849 8435 11883
rect 8435 11849 8444 11883
rect 8392 11840 8444 11849
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 1492 11636 1544 11688
rect 1860 11636 1912 11688
rect 2136 11704 2188 11756
rect 2320 11704 2372 11756
rect 2872 11704 2924 11756
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 5632 11704 5684 11756
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 2412 11568 2464 11620
rect 7196 11568 7248 11620
rect 10416 11611 10468 11620
rect 10416 11577 10425 11611
rect 10425 11577 10459 11611
rect 10459 11577 10468 11611
rect 10416 11568 10468 11577
rect 1768 11500 1820 11552
rect 2136 11500 2188 11552
rect 7104 11500 7156 11552
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 9312 11500 9364 11552
rect 10140 11500 10192 11552
rect 11152 11500 11204 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1676 11296 1728 11348
rect 5632 11339 5684 11348
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 9772 11296 9824 11348
rect 10600 11296 10652 11348
rect 1860 11228 1912 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 7840 11228 7892 11280
rect 9312 11228 9364 11280
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 7012 11092 7064 11144
rect 7380 11092 7432 11144
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 8668 11092 8720 11144
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9496 11092 9548 11144
rect 9680 11024 9732 11076
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 7564 10956 7616 10965
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 1768 10752 1820 10804
rect 2228 10752 2280 10804
rect 5264 10752 5316 10804
rect 7196 10752 7248 10804
rect 8024 10752 8076 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 1768 10616 1820 10668
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 2688 10616 2740 10668
rect 4252 10684 4304 10736
rect 3884 10616 3936 10668
rect 2412 10548 2464 10600
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 7840 10616 7892 10668
rect 8668 10616 8720 10668
rect 9680 10752 9732 10804
rect 10692 10752 10744 10804
rect 9772 10727 9824 10736
rect 9772 10693 9806 10727
rect 9806 10693 9824 10727
rect 9772 10684 9824 10693
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 8300 10548 8352 10600
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 7196 10480 7248 10532
rect 8116 10480 8168 10532
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 1584 10208 1636 10260
rect 3884 10208 3936 10260
rect 1308 10140 1360 10192
rect 1584 10004 1636 10056
rect 2504 10072 2556 10124
rect 2688 10072 2740 10124
rect 6460 10072 6512 10124
rect 6828 10072 6880 10124
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 7564 10004 7616 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8300 10047 8352 10056
rect 8300 10013 8317 10047
rect 8317 10013 8351 10047
rect 8351 10013 8352 10047
rect 8300 10004 8352 10013
rect 9128 9936 9180 9988
rect 1768 9868 1820 9920
rect 7564 9868 7616 9920
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 11152 9868 11204 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 7748 9596 7800 9648
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 6828 9528 6880 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10140 9596 10192 9648
rect 10048 9528 10100 9580
rect 9588 9460 9640 9512
rect 7012 9392 7064 9444
rect 9496 9392 9548 9444
rect 1308 9324 1360 9376
rect 9220 9324 9272 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 10692 9120 10744 9172
rect 1768 9052 1820 9104
rect 1308 8916 1360 8968
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 2320 8916 2372 8968
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 9220 9027 9272 9036
rect 9220 8993 9229 9027
rect 9229 8993 9263 9027
rect 9263 8993 9272 9027
rect 9220 8984 9272 8993
rect 9496 8984 9548 9036
rect 4160 8916 4212 8968
rect 7012 8916 7064 8968
rect 7564 8959 7616 8968
rect 7564 8925 7598 8959
rect 7598 8925 7616 8959
rect 7564 8916 7616 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 2228 8823 2280 8832
rect 2228 8789 2237 8823
rect 2237 8789 2271 8823
rect 2271 8789 2280 8823
rect 2228 8780 2280 8789
rect 10968 8823 11020 8832
rect 10968 8789 10977 8823
rect 10977 8789 11011 8823
rect 11011 8789 11020 8823
rect 10968 8780 11020 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2412 8576 2464 8628
rect 2688 8576 2740 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 9128 8508 9180 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 2780 8440 2832 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 10048 8551 10100 8560
rect 10048 8517 10057 8551
rect 10057 8517 10091 8551
rect 10091 8517 10100 8551
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 10048 8508 10100 8517
rect 10140 8440 10192 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 2320 8304 2372 8356
rect 9312 8372 9364 8424
rect 9036 8304 9088 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 2780 7964 2832 8016
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 10508 7828 10560 7880
rect 848 7692 900 7744
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1676 7488 1728 7540
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 11060 7488 11112 7540
rect 1308 7352 1360 7404
rect 3240 7352 3292 7404
rect 4160 7352 4212 7404
rect 9496 7420 9548 7472
rect 9220 7352 9272 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 10508 7259 10560 7268
rect 10508 7225 10517 7259
rect 10517 7225 10551 7259
rect 10551 7225 10560 7259
rect 10508 7216 10560 7225
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 11060 7148 11112 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2320 6944 2372 6996
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 3240 6919 3292 6928
rect 3240 6885 3249 6919
rect 3249 6885 3283 6919
rect 3283 6885 3292 6919
rect 3240 6876 3292 6885
rect 2688 6808 2740 6860
rect 8760 6808 8812 6860
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 9312 6740 9364 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 1584 6672 1636 6724
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 2872 6400 2924 6452
rect 9220 6400 9272 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 1308 6264 1360 6316
rect 1676 6332 1728 6384
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 8208 6264 8260 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 10232 6264 10284 6316
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 8668 6060 8720 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1308 5856 1360 5908
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 9312 5856 9364 5908
rect 10232 5899 10284 5908
rect 10232 5865 10241 5899
rect 10241 5865 10275 5899
rect 10275 5865 10284 5899
rect 10232 5856 10284 5865
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 8576 5720 8628 5772
rect 1400 5652 1452 5661
rect 1768 5516 1820 5568
rect 8576 5627 8628 5636
rect 8576 5593 8585 5627
rect 8585 5593 8619 5627
rect 8619 5593 8628 5627
rect 8576 5584 8628 5593
rect 8760 5627 8812 5636
rect 8760 5593 8769 5627
rect 8769 5593 8803 5627
rect 8803 5593 8812 5627
rect 8760 5584 8812 5593
rect 10416 5652 10468 5704
rect 11152 5652 11204 5704
rect 8668 5516 8720 5568
rect 9404 5516 9456 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2688 5355 2740 5364
rect 2688 5321 2697 5355
rect 2697 5321 2731 5355
rect 2731 5321 2740 5355
rect 2688 5312 2740 5321
rect 1768 5287 1820 5296
rect 1768 5253 1777 5287
rect 1777 5253 1811 5287
rect 1811 5253 1820 5287
rect 1768 5244 1820 5253
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 6920 5244 6972 5296
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 9680 5176 9732 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 1860 5108 1912 5160
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 6736 5108 6788 5160
rect 9588 5108 9640 5160
rect 4804 4972 4856 5024
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2964 4768 3016 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 1308 4564 1360 4616
rect 1860 4564 1912 4616
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 6736 4539 6788 4548
rect 6736 4505 6745 4539
rect 6745 4505 6779 4539
rect 6779 4505 6788 4539
rect 6736 4496 6788 4505
rect 9864 4539 9916 4548
rect 9864 4505 9898 4539
rect 9898 4505 9916 4539
rect 9864 4496 9916 4505
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 10140 4224 10192 4276
rect 1216 4088 1268 4140
rect 4620 4088 4672 4140
rect 1584 4020 1636 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 2688 4063 2740 4072
rect 2688 4029 2697 4063
rect 2697 4029 2731 4063
rect 2731 4029 2740 4063
rect 2688 4020 2740 4029
rect 4068 4020 4120 4072
rect 3056 3952 3108 4004
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 10324 4156 10376 4208
rect 10784 4088 10836 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 1676 3884 1728 3936
rect 5264 3884 5316 3936
rect 7564 3884 7616 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2688 3680 2740 3732
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 10140 3680 10192 3732
rect 10968 3680 11020 3732
rect 2596 3612 2648 3664
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 10784 3655 10836 3664
rect 10784 3621 10793 3655
rect 10793 3621 10827 3655
rect 10827 3621 10836 3655
rect 10784 3612 10836 3621
rect 3148 3544 3200 3596
rect 3516 3544 3568 3596
rect 1676 3476 1728 3485
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4160 3408 4212 3460
rect 6736 3544 6788 3596
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 5264 3451 5316 3460
rect 5264 3417 5298 3451
rect 5298 3417 5316 3451
rect 5264 3408 5316 3417
rect 5724 3408 5776 3460
rect 7564 3476 7616 3528
rect 8760 3476 8812 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 6920 3408 6972 3460
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 4620 3340 4672 3392
rect 6368 3383 6420 3392
rect 6368 3349 6377 3383
rect 6377 3349 6411 3383
rect 6411 3349 6420 3383
rect 6368 3340 6420 3349
rect 6552 3383 6604 3392
rect 6552 3349 6561 3383
rect 6561 3349 6595 3383
rect 6595 3349 6604 3383
rect 6552 3340 6604 3349
rect 8484 3340 8536 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1492 3136 1544 3188
rect 4068 3136 4120 3188
rect 6460 3136 6512 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 2780 3068 2832 3120
rect 8024 3068 8076 3120
rect 1308 3000 1360 3052
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5540 3000 5592 3052
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 8392 3000 8444 3052
rect 9496 3068 9548 3120
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 7196 2864 7248 2916
rect 4160 2796 4212 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 4620 2592 4672 2644
rect 4712 2592 4764 2644
rect 5540 2592 5592 2644
rect 8024 2592 8076 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 8392 2592 8444 2644
rect 9680 2592 9732 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 11060 2592 11112 2644
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 2872 2320 2924 2372
rect 4804 2388 4856 2440
rect 6368 2388 6420 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8208 2524 8260 2576
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 5264 2252 5316 2304
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 8392 2252 8444 2304
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9036 2252 9088 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5170 13767 5226 14567
rect 5814 13767 5870 14567
rect 6458 13767 6514 14567
rect 7102 13767 7158 14567
rect 7746 13767 7802 14567
rect 8390 13767 8446 14567
rect 9034 13767 9090 14567
rect 2870 13016 2926 13025
rect 2870 12951 2926 12960
rect 1030 12336 1086 12345
rect 1030 12271 1086 12280
rect 1044 11898 1072 12271
rect 2884 11898 2912 12951
rect 5184 12186 5212 13767
rect 5184 12158 5304 12186
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11898 5304 12158
rect 5828 11898 5856 13767
rect 6472 11898 6500 13767
rect 7116 11898 7144 13767
rect 7760 11898 7788 13767
rect 8404 11898 8432 13767
rect 9048 11898 9076 13767
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 1032 11892 1084 11898
rect 1032 11834 1084 11840
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 2884 11762 2912 11834
rect 10244 11762 10272 12951
rect 11058 12336 11114 12345
rect 11058 12271 11114 12280
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 11218 1532 11630
rect 1688 11354 1716 11698
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1780 10810 1808 11494
rect 1872 11286 1900 11630
rect 2148 11558 2176 11698
rect 2332 11665 2360 11698
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 2148 10985 2176 11494
rect 2424 11150 2452 11562
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 2134 10976 2190 10985
rect 2134 10911 2190 10920
rect 2240 10810 2268 11086
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1780 10674 1808 10746
rect 4264 10742 4292 11086
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10810 5304 11698
rect 5644 11354 5672 11698
rect 10414 11656 10470 11665
rect 7196 11620 7248 11626
rect 10414 11591 10416 11600
rect 7196 11562 7248 11568
rect 10468 11591 10470 11600
rect 10416 11562 10468 11568
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 1306 10296 1362 10305
rect 1596 10266 1624 10610
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 1306 10231 1362 10240
rect 1584 10260 1636 10266
rect 1320 10198 1348 10231
rect 1584 10202 1636 10208
rect 1308 10192 1360 10198
rect 1308 10134 1360 10140
rect 2424 10062 2452 10542
rect 2516 10130 2544 10610
rect 2700 10130 2728 10610
rect 3896 10266 3924 10610
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 6840 10130 6868 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 1596 9654 1624 9998
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1584 9648 1636 9654
rect 1582 9616 1584 9625
rect 1636 9616 1638 9625
rect 1582 9551 1638 9560
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1320 8974 1348 9318
rect 1780 9110 1808 9862
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1780 8974 1808 9046
rect 1308 8968 1360 8974
rect 1306 8936 1308 8945
rect 1768 8968 1820 8974
rect 1360 8936 1362 8945
rect 1768 8910 1820 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 1306 8871 1362 8880
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 2240 7886 2268 8774
rect 2332 8498 2360 8910
rect 2424 8634 2452 8910
rect 2700 8634 2728 10066
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 6472 9586 6500 10066
rect 6840 9586 6868 10066
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 4172 8498 4200 8910
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 7954 2360 8298
rect 2792 8022 2820 8434
rect 4172 8378 4200 8434
rect 4080 8350 4200 8378
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 4080 7970 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2320 7948 2372 7954
rect 4080 7942 4200 7970
rect 2320 7890 2372 7896
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1688 7546 1716 7822
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 6905 1348 7346
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6914 1624 7142
rect 2332 7002 2360 7890
rect 4172 7410 4200 7942
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 6932 7546 6960 9522
rect 7024 9450 7052 11086
rect 7116 10690 7144 11494
rect 7208 11218 7236 11562
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7208 10810 7236 11154
rect 7392 11150 7420 11494
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7852 11150 7880 11222
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7116 10674 7236 10690
rect 7392 10674 7420 11086
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7116 10668 7248 10674
rect 7116 10662 7196 10668
rect 7196 10610 7248 10616
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7208 10538 7236 10610
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7576 10062 7604 10950
rect 7852 10674 7880 11086
rect 8036 10810 8064 11086
rect 8312 10810 8340 11154
rect 8680 11150 8708 11494
rect 9324 11286 9352 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9324 11150 9352 11222
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8680 10674 8708 11086
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9508 10606 9536 11086
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10810 9720 11018
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 10742 9812 11290
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 8974 7052 9386
rect 7576 8974 7604 9862
rect 7760 9654 7788 10066
rect 8128 10062 8156 10474
rect 8312 10062 8340 10542
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 9140 8974 9168 9930
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9042 9260 9318
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8566 9168 8910
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9324 8430 9352 9522
rect 9508 9450 9536 10542
rect 10152 9654 10180 11494
rect 10612 11354 10640 11698
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10704 10810 10732 11698
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10598 10296 10654 10305
rect 10598 10231 10654 10240
rect 10612 10062 10640 10231
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9042 9536 9386
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 3252 6934 3280 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3240 6928 3292 6934
rect 1306 6896 1362 6905
rect 1596 6886 1716 6914
rect 1306 6831 1362 6840
rect 1688 6798 1716 6886
rect 3240 6870 3292 6876
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1596 6458 1624 6666
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1688 6390 1716 6734
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6458 1992 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 2332 6322 2360 6734
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1320 6225 1348 6258
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1320 5914 1348 6151
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1768 5568 1820 5574
rect 1398 5536 1454 5545
rect 1768 5510 1820 5516
rect 1398 5471 1454 5480
rect 1780 5302 1808 5510
rect 2700 5370 2728 6802
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2884 6458 2912 6734
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 6932 5302 6960 7482
rect 9048 6866 9076 8298
rect 9508 7478 9536 8978
rect 9600 8634 9628 9454
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 10060 8566 10088 9522
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10152 8498 10180 9590
rect 10704 9178 10732 9998
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10796 8634 10824 8871
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10980 8498 11008 8774
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10612 8265 10640 8434
rect 10598 8256 10654 8265
rect 10598 8191 10654 8200
rect 10612 8090 10640 8191
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8772 6322 8800 6802
rect 9232 6458 9260 7346
rect 10520 7274 10548 7822
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7585 10916 7686
rect 10874 7576 10930 7585
rect 11072 7546 11100 12271
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 10985 11192 11494
rect 11150 10976 11206 10985
rect 11150 10911 11206 10920
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9625 11192 9862
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 10874 7511 10930 7520
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10980 7002 11008 7346
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11072 6905 11100 7142
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9324 6458 9352 6734
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8220 5914 8248 6258
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8588 5778 8616 6054
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5658 8708 6054
rect 9324 5914 9352 6258
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8588 5642 8708 5658
rect 8576 5636 8708 5642
rect 8628 5630 8708 5636
rect 8760 5636 8812 5642
rect 8576 5578 8628 5584
rect 8760 5578 8812 5584
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1306 4856 1362 4865
rect 1596 4826 1624 5170
rect 1306 4791 1362 4800
rect 1584 4820 1636 4826
rect 1320 4622 1348 4791
rect 1584 4762 1636 4768
rect 1780 4706 1808 5238
rect 8588 5234 8616 5578
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5370 8708 5510
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8772 5234 8800 5578
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1872 4826 1900 5102
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1780 4678 1900 4706
rect 1872 4622 1900 4678
rect 2424 4622 2452 5170
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2884 4282 2912 5102
rect 2976 4826 3004 5170
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 1214 4176 1270 4185
rect 1214 4111 1216 4120
rect 1268 4111 1270 4120
rect 1216 4082 1268 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 1596 3738 1624 4014
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1688 3534 1716 3878
rect 2608 3670 2636 4014
rect 2700 3738 2728 4014
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 3068 3534 3096 3946
rect 3528 3602 3556 5102
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3618 4108 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3738 4660 4082
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3516 3596 3568 3602
rect 4080 3590 4200 3618
rect 3516 3538 3568 3544
rect 1492 3528 1544 3534
rect 1306 3496 1362 3505
rect 1492 3470 1544 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 1306 3431 1362 3440
rect 1320 3058 1348 3431
rect 1504 3194 1532 3470
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 2792 3126 2820 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3160 3058 3188 3538
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3194 4108 3470
rect 4172 3466 4200 3590
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2884 2378 2912 2994
rect 3068 2650 3096 2994
rect 4172 2854 4200 3402
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 3334
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4724 2650 4752 2994
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4816 2446 4844 4966
rect 6748 4554 6776 5102
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3466 5304 3878
rect 6748 3602 6776 4490
rect 9416 4078 9444 5510
rect 9600 5166 9628 6734
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10244 5914 10272 6258
rect 10980 6225 11008 6258
rect 10966 6216 11022 6225
rect 10966 6151 11022 6160
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4690 9628 5102
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7576 3534 7604 3878
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5552 2650 5580 2994
rect 5736 2990 5764 3402
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 6380 2446 6408 3334
rect 6472 3194 6500 3470
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6564 3058 6592 3334
rect 6932 3194 6960 3402
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7576 3058 7604 3470
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8036 2990 8064 3062
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7208 2446 7236 2858
rect 8036 2650 8064 2926
rect 8312 2650 8340 2994
rect 8404 2650 8432 2994
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8208 2576 8260 2582
rect 8404 2530 8432 2586
rect 8260 2524 8432 2530
rect 8208 2518 8432 2524
rect 8220 2502 8432 2518
rect 8496 2446 8524 3334
rect 8772 3194 8800 3470
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9508 3126 9536 3334
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9600 3058 9628 4626
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9692 2650 9720 5170
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 4282 9904 4490
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10152 4146 10180 4218
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3738 10180 4082
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10336 3534 10364 4150
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10428 2650 10456 5646
rect 11164 5545 11192 5646
rect 11150 5536 11206 5545
rect 11150 5471 11206 5480
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4865 10824 4966
rect 10782 4856 10838 4865
rect 10980 4826 11008 5170
rect 10782 4791 10838 4800
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10966 4176 11022 4185
rect 10784 4140 10836 4146
rect 10966 4111 10968 4120
rect 10784 4082 10836 4088
rect 11020 4111 11022 4120
rect 10968 4082 11020 4088
rect 10796 3670 10824 4082
rect 10980 3738 11008 4082
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10968 3528 11020 3534
rect 10966 3496 10968 3505
rect 11020 3496 11022 3505
rect 10966 3431 11022 3440
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11058 2816 11114 2825
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10980 2446 11008 2790
rect 11058 2751 11114 2760
rect 11072 2650 11100 2751
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 3252 800 3280 2382
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 3896 800 3924 2246
rect 4540 800 4568 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1170 5304 2246
rect 5184 1142 5304 1170
rect 5184 800 5212 1142
rect 5828 800 5856 2246
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 9048 800 9076 2246
rect 10336 2145 10364 2382
rect 10322 2136 10378 2145
rect 10322 2071 10378 2080
rect 10612 1465 10640 2382
rect 10598 1456 10654 1465
rect 10598 1391 10654 1400
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
<< via2 >>
rect 2870 12960 2926 13016
rect 1030 12280 1086 12336
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 10230 12960 10286 13016
rect 11058 12280 11114 12336
rect 2318 11600 2374 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 2134 10920 2190 10976
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 10414 11620 10470 11656
rect 10414 11600 10416 11620
rect 10416 11600 10468 11620
rect 10468 11600 10470 11620
rect 1306 10240 1362 10296
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1582 9596 1584 9616
rect 1584 9596 1636 9616
rect 1636 9596 1638 9616
rect 1582 9560 1638 9596
rect 1306 8916 1308 8936
rect 1308 8916 1360 8936
rect 1360 8916 1362 8936
rect 1306 8880 1362 8916
rect 1490 8200 1546 8256
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 10598 10240 10654 10296
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1306 6840 1362 6896
rect 1306 6160 1362 6216
rect 1398 5480 1454 5536
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 10782 8880 10838 8936
rect 10598 8200 10654 8256
rect 10874 7520 10930 7576
rect 11150 10920 11206 10976
rect 11150 9560 11206 9616
rect 11058 6840 11114 6896
rect 1306 4800 1362 4856
rect 1214 4140 1270 4176
rect 1214 4120 1216 4140
rect 1216 4120 1268 4140
rect 1268 4120 1270 4140
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1306 3440 1362 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 10966 6160 11022 6216
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 11150 5480 11206 5536
rect 10782 4800 10838 4856
rect 10966 4140 11022 4176
rect 10966 4120 10968 4140
rect 10968 4120 11020 4140
rect 11020 4120 11022 4140
rect 10966 3476 10968 3496
rect 10968 3476 11020 3496
rect 11020 3476 11022 3496
rect 10966 3440 11022 3476
rect 11058 2760 11114 2816
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 10322 2080 10378 2136
rect 10598 1400 10654 1456
<< metal3 >>
rect 0 13018 800 13048
rect 2865 13018 2931 13021
rect 0 13016 2931 13018
rect 0 12960 2870 13016
rect 2926 12960 2931 13016
rect 0 12958 2931 12960
rect 0 12928 800 12958
rect 2865 12955 2931 12958
rect 10225 13018 10291 13021
rect 11623 13018 12423 13048
rect 10225 13016 12423 13018
rect 10225 12960 10230 13016
rect 10286 12960 12423 13016
rect 10225 12958 12423 12960
rect 10225 12955 10291 12958
rect 11623 12928 12423 12958
rect 0 12338 800 12368
rect 1025 12338 1091 12341
rect 0 12336 1091 12338
rect 0 12280 1030 12336
rect 1086 12280 1091 12336
rect 0 12278 1091 12280
rect 0 12248 800 12278
rect 1025 12275 1091 12278
rect 11053 12338 11119 12341
rect 11623 12338 12423 12368
rect 11053 12336 12423 12338
rect 11053 12280 11058 12336
rect 11114 12280 12423 12336
rect 11053 12278 12423 12280
rect 11053 12275 11119 12278
rect 11623 12248 12423 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 2313 11658 2379 11661
rect 0 11656 2379 11658
rect 0 11600 2318 11656
rect 2374 11600 2379 11656
rect 0 11598 2379 11600
rect 0 11568 800 11598
rect 2313 11595 2379 11598
rect 10409 11658 10475 11661
rect 11623 11658 12423 11688
rect 10409 11656 12423 11658
rect 10409 11600 10414 11656
rect 10470 11600 12423 11656
rect 10409 11598 12423 11600
rect 10409 11595 10475 11598
rect 11623 11568 12423 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 0 10978 800 11008
rect 2129 10978 2195 10981
rect 0 10976 2195 10978
rect 0 10920 2134 10976
rect 2190 10920 2195 10976
rect 0 10918 2195 10920
rect 0 10888 800 10918
rect 2129 10915 2195 10918
rect 11145 10978 11211 10981
rect 11623 10978 12423 11008
rect 11145 10976 12423 10978
rect 11145 10920 11150 10976
rect 11206 10920 12423 10976
rect 11145 10918 12423 10920
rect 11145 10915 11211 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 11623 10888 12423 10918
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 10593 10298 10659 10301
rect 11623 10298 12423 10328
rect 10593 10296 12423 10298
rect 10593 10240 10598 10296
rect 10654 10240 12423 10296
rect 10593 10238 12423 10240
rect 10593 10235 10659 10238
rect 11623 10208 12423 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 11145 9618 11211 9621
rect 11623 9618 12423 9648
rect 11145 9616 12423 9618
rect 11145 9560 11150 9616
rect 11206 9560 12423 9616
rect 11145 9558 12423 9560
rect 11145 9555 11211 9558
rect 11623 9528 12423 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 10777 8938 10843 8941
rect 11623 8938 12423 8968
rect 10777 8936 12423 8938
rect 10777 8880 10782 8936
rect 10838 8880 12423 8936
rect 10777 8878 12423 8880
rect 10777 8875 10843 8878
rect 11623 8848 12423 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 10593 8258 10659 8261
rect 11623 8258 12423 8288
rect 10593 8256 12423 8258
rect 10593 8200 10598 8256
rect 10654 8200 12423 8256
rect 10593 8198 12423 8200
rect 10593 8195 10659 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 11623 8168 12423 8198
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 10869 7578 10935 7581
rect 11623 7578 12423 7608
rect 10869 7576 12423 7578
rect 10869 7520 10874 7576
rect 10930 7520 12423 7576
rect 10869 7518 12423 7520
rect 0 7488 800 7518
rect 10869 7515 10935 7518
rect 11623 7488 12423 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 800 6838
rect 1301 6835 1367 6838
rect 11053 6898 11119 6901
rect 11623 6898 12423 6928
rect 11053 6896 12423 6898
rect 11053 6840 11058 6896
rect 11114 6840 12423 6896
rect 11053 6838 12423 6840
rect 11053 6835 11119 6838
rect 11623 6808 12423 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 10961 6218 11027 6221
rect 11623 6218 12423 6248
rect 10961 6216 12423 6218
rect 10961 6160 10966 6216
rect 11022 6160 12423 6216
rect 10961 6158 12423 6160
rect 10961 6155 11027 6158
rect 11623 6128 12423 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 11145 5538 11211 5541
rect 11623 5538 12423 5568
rect 11145 5536 12423 5538
rect 11145 5480 11150 5536
rect 11206 5480 12423 5536
rect 11145 5478 12423 5480
rect 11145 5475 11211 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 11623 5448 12423 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 10777 4858 10843 4861
rect 11623 4858 12423 4888
rect 10777 4856 12423 4858
rect 10777 4800 10782 4856
rect 10838 4800 12423 4856
rect 10777 4798 12423 4800
rect 10777 4795 10843 4798
rect 11623 4768 12423 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1209 4178 1275 4181
rect 0 4176 1275 4178
rect 0 4120 1214 4176
rect 1270 4120 1275 4176
rect 0 4118 1275 4120
rect 0 4088 800 4118
rect 1209 4115 1275 4118
rect 10961 4178 11027 4181
rect 11623 4178 12423 4208
rect 10961 4176 12423 4178
rect 10961 4120 10966 4176
rect 11022 4120 12423 4176
rect 10961 4118 12423 4120
rect 10961 4115 11027 4118
rect 11623 4088 12423 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 0 3498 800 3528
rect 1301 3498 1367 3501
rect 0 3496 1367 3498
rect 0 3440 1306 3496
rect 1362 3440 1367 3496
rect 0 3438 1367 3440
rect 0 3408 800 3438
rect 1301 3435 1367 3438
rect 10961 3498 11027 3501
rect 11623 3498 12423 3528
rect 10961 3496 12423 3498
rect 10961 3440 10966 3496
rect 11022 3440 12423 3496
rect 10961 3438 12423 3440
rect 10961 3435 11027 3438
rect 11623 3408 12423 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 11053 2818 11119 2821
rect 11623 2818 12423 2848
rect 11053 2816 12423 2818
rect 11053 2760 11058 2816
rect 11114 2760 12423 2816
rect 11053 2758 12423 2760
rect 11053 2755 11119 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 11623 2728 12423 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 10317 2138 10383 2141
rect 11623 2138 12423 2168
rect 10317 2136 12423 2138
rect 10317 2080 10322 2136
rect 10378 2080 12423 2136
rect 10317 2078 12423 2080
rect 10317 2075 10383 2078
rect 11623 2048 12423 2078
rect 10593 1458 10659 1461
rect 11623 1458 12423 1488
rect 10593 1456 12423 1458
rect 10593 1400 10598 1456
rect 10654 1400 12423 1456
rect 10593 1398 12423 1400
rect 10593 1395 10659 1398
rect 11623 1368 12423 1398
<< via3 >>
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect -2966 16006 -2346 16038
rect -2966 15770 -2934 16006
rect -2698 15770 -2614 16006
rect -2378 15770 -2346 16006
rect -2966 15686 -2346 15770
rect -2966 15450 -2934 15686
rect -2698 15450 -2614 15686
rect -2378 15450 -2346 15686
rect -2966 6284 -2346 15450
rect -2966 6048 -2934 6284
rect -2698 6048 -2614 6284
rect -2378 6048 -2346 6284
rect -2966 -1306 -2346 6048
rect -2006 15046 -1386 15078
rect -2006 14810 -1974 15046
rect -1738 14810 -1654 15046
rect -1418 14810 -1386 15046
rect -2006 14726 -1386 14810
rect -2006 14490 -1974 14726
rect -1738 14490 -1654 14726
rect -1418 14490 -1386 14726
rect -2006 5624 -1386 14490
rect -2006 5388 -1974 5624
rect -1738 5388 -1654 5624
rect -1418 5388 -1386 5624
rect -2006 -346 -1386 5388
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 4208 15046 4528 16038
rect 4208 14810 4250 15046
rect 4486 14810 4528 15046
rect 4208 14726 4528 14810
rect 4208 14490 4250 14726
rect 4486 14490 4528 14726
rect 4208 11456 4528 14490
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 -346 4528 2688
rect 4208 -582 4250 -346
rect 4486 -582 4528 -346
rect 4208 -666 4528 -582
rect 4208 -902 4250 -666
rect 4486 -902 4528 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 4208 -1894 4528 -902
rect 4868 16006 5188 16038
rect 4868 15770 4910 16006
rect 5146 15770 5188 16006
rect 4868 15686 5188 15770
rect 4868 15450 4910 15686
rect 5146 15450 5188 15686
rect 4868 12000 5188 15450
rect 14766 16006 15386 16038
rect 14766 15770 14798 16006
rect 15034 15770 15118 16006
rect 15354 15770 15386 16006
rect 14766 15686 15386 15770
rect 14766 15450 14798 15686
rect 15034 15450 15118 15686
rect 15354 15450 15386 15686
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 -1306 5188 2144
rect 13806 15046 14426 15078
rect 13806 14810 13838 15046
rect 14074 14810 14158 15046
rect 14394 14810 14426 15046
rect 13806 14726 14426 14810
rect 13806 14490 13838 14726
rect 14074 14490 14158 14726
rect 14394 14490 14426 14726
rect 13806 5624 14426 14490
rect 13806 5388 13838 5624
rect 14074 5388 14158 5624
rect 14394 5388 14426 5624
rect 13806 -346 14426 5388
rect 13806 -582 13838 -346
rect 14074 -582 14158 -346
rect 14394 -582 14426 -346
rect 13806 -666 14426 -582
rect 13806 -902 13838 -666
rect 14074 -902 14158 -666
rect 14394 -902 14426 -666
rect 13806 -934 14426 -902
rect 14766 6284 15386 15450
rect 14766 6048 14798 6284
rect 15034 6048 15118 6284
rect 15354 6048 15386 6284
rect 4868 -1542 4910 -1306
rect 5146 -1542 5188 -1306
rect 4868 -1626 5188 -1542
rect 4868 -1862 4910 -1626
rect 5146 -1862 5188 -1626
rect 4868 -1894 5188 -1862
rect 14766 -1306 15386 6048
rect 14766 -1542 14798 -1306
rect 15034 -1542 15118 -1306
rect 15354 -1542 15386 -1306
rect 14766 -1626 15386 -1542
rect 14766 -1862 14798 -1626
rect 15034 -1862 15118 -1626
rect 15354 -1862 15386 -1626
rect 14766 -1894 15386 -1862
<< via4 >>
rect -2934 15770 -2698 16006
rect -2614 15770 -2378 16006
rect -2934 15450 -2698 15686
rect -2614 15450 -2378 15686
rect -2934 6048 -2698 6284
rect -2614 6048 -2378 6284
rect -1974 14810 -1738 15046
rect -1654 14810 -1418 15046
rect -1974 14490 -1738 14726
rect -1654 14490 -1418 14726
rect -1974 5388 -1738 5624
rect -1654 5388 -1418 5624
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 4250 14810 4486 15046
rect 4250 14490 4486 14726
rect 4250 5388 4486 5624
rect 4250 -582 4486 -346
rect 4250 -902 4486 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4910 15770 5146 16006
rect 4910 15450 5146 15686
rect 14798 15770 15034 16006
rect 15118 15770 15354 16006
rect 14798 15450 15034 15686
rect 15118 15450 15354 15686
rect 4910 6048 5146 6284
rect 13838 14810 14074 15046
rect 14158 14810 14394 15046
rect 13838 14490 14074 14726
rect 14158 14490 14394 14726
rect 13838 5388 14074 5624
rect 14158 5388 14394 5624
rect 13838 -582 14074 -346
rect 14158 -582 14394 -346
rect 13838 -902 14074 -666
rect 14158 -902 14394 -666
rect 14798 6048 15034 6284
rect 15118 6048 15354 6284
rect 4910 -1542 5146 -1306
rect 4910 -1862 5146 -1626
rect 14798 -1542 15034 -1306
rect 15118 -1542 15354 -1306
rect 14798 -1862 15034 -1626
rect 15118 -1862 15354 -1626
<< metal5 >>
rect -2966 16006 15386 16038
rect -2966 15770 -2934 16006
rect -2698 15770 -2614 16006
rect -2378 15770 4910 16006
rect 5146 15770 14798 16006
rect 15034 15770 15118 16006
rect 15354 15770 15386 16006
rect -2966 15686 15386 15770
rect -2966 15450 -2934 15686
rect -2698 15450 -2614 15686
rect -2378 15450 4910 15686
rect 5146 15450 14798 15686
rect 15034 15450 15118 15686
rect 15354 15450 15386 15686
rect -2966 15418 15386 15450
rect -2006 15046 14426 15078
rect -2006 14810 -1974 15046
rect -1738 14810 -1654 15046
rect -1418 14810 4250 15046
rect 4486 14810 13838 15046
rect 14074 14810 14158 15046
rect 14394 14810 14426 15046
rect -2006 14726 14426 14810
rect -2006 14490 -1974 14726
rect -1738 14490 -1654 14726
rect -1418 14490 4250 14726
rect 4486 14490 13838 14726
rect 14074 14490 14158 14726
rect 14394 14490 14426 14726
rect -2006 14458 14426 14490
rect -2966 6284 15386 6326
rect -2966 6048 -2934 6284
rect -2698 6048 -2614 6284
rect -2378 6048 4910 6284
rect 5146 6048 14798 6284
rect 15034 6048 15118 6284
rect 15354 6048 15386 6284
rect -2966 6006 15386 6048
rect -2966 5624 15386 5666
rect -2966 5388 -1974 5624
rect -1738 5388 -1654 5624
rect -1418 5388 4250 5624
rect 4486 5388 13838 5624
rect 14074 5388 14158 5624
rect 14394 5388 15386 5624
rect -2966 5346 15386 5388
rect -2006 -346 14426 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 4250 -346
rect 4486 -582 13838 -346
rect 14074 -582 14158 -346
rect 14394 -582 14426 -346
rect -2006 -666 14426 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 4250 -666
rect 4486 -902 13838 -666
rect 14074 -902 14158 -666
rect 14394 -902 14426 -666
rect -2006 -934 14426 -902
rect -2966 -1306 15386 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 4910 -1306
rect 5146 -1542 14798 -1306
rect 15034 -1542 15118 -1306
rect 15354 -1542 15386 -1306
rect -2966 -1626 15386 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 4910 -1626
rect 5146 -1862 14798 -1626
rect 15034 -1862 15118 -1626
rect 15354 -1862 15386 -1626
rect -2966 -1894 15386 -1862
use sky130_fd_sc_hd__and2_1  _060_
timestamp -3599
transform 1 0 7268 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _061_
timestamp -3599
transform 1 0 6900 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _062_
timestamp -3599
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _063_
timestamp -3599
transform 1 0 8188 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _064_
timestamp -3599
transform 1 0 7544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _065_
timestamp -3599
transform -1 0 7268 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _066_
timestamp -3599
transform 1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _067_
timestamp -3599
transform 1 0 6440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _068_
timestamp -3599
transform -1 0 8096 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _069_
timestamp -3599
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _070_
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _071_
timestamp -3599
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _072_
timestamp -3599
transform -1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _073_
timestamp -3599
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _074_
timestamp -3599
transform -1 0 10120 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _075_
timestamp -3599
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _076_
timestamp -3599
transform -1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _077_
timestamp -3599
transform -1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _078_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _079_
timestamp -3599
transform -1 0 8832 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _080_
timestamp -3599
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _081_
timestamp -3599
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _082_
timestamp -3599
transform -1 0 9292 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _083_
timestamp -3599
transform 1 0 7912 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp -3599
transform -1 0 10672 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _085_
timestamp -3599
transform 1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _086_
timestamp -3599
transform -1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _087_
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _088_
timestamp -3599
transform 1 0 9292 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _089_
timestamp -3599
transform -1 0 8556 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp -3599
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _091_
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _092_
timestamp -3599
transform -1 0 9292 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _093_
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _094_
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _095_
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _096_
timestamp -3599
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _097_
timestamp -3599
transform -1 0 8096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _098_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _099_
timestamp -3599
transform -1 0 3128 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _101_
timestamp -3599
transform -1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _102_
timestamp -3599
transform -1 0 6164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _103_
timestamp -3599
transform 1 0 4048 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp -3599
transform 1 0 1748 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _105_
timestamp -3599
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _106_
timestamp -3599
transform -1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _107_
timestamp -3599
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _108_
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _109_
timestamp -3599
transform 1 0 1564 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _110_
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _111_
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _112_
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _113_
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _114_
timestamp -3599
transform 1 0 1472 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _115_
timestamp -3599
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _116_
timestamp -3599
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _117_
timestamp -3599
transform 1 0 2024 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _118_
timestamp -3599
transform 1 0 2668 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _119_
timestamp -3599
transform 1 0 1748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _120_
timestamp -3599
transform -1 0 2760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp -3599
transform -1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _122_
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _123_
timestamp -3599
transform 1 0 2024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _124_
timestamp -3599
transform 1 0 1656 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _125_
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _126_
timestamp -3599
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _127_
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _128_
timestamp -3599
transform 1 0 2668 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _129_
timestamp -3599
transform 1 0 1472 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _130_
timestamp -3599
transform -1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp -3599
transform -1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _132_
timestamp -3599
transform 1 0 2116 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _133_
timestamp -3599
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _134_
timestamp -3599
transform 1 0 2852 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _135_
timestamp -3599
transform -1 0 9384 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _136_
timestamp -3599
transform 1 0 8740 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _137_
timestamp -3599
transform 1 0 9568 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp -3599
transform 1 0 9476 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp -3599
transform 1 0 7268 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp -3599
transform 1 0 9568 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp -3599
transform 1 0 9568 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp -3599
transform 1 0 9108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _143_
timestamp -3599
transform 1 0 9568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _144_
timestamp -3599
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _145_
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _146_
timestamp -3599
transform 1 0 4968 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _147_
timestamp -3599
transform 1 0 3128 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _148_
timestamp -3599
transform 1 0 3496 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _149_
timestamp -3599
transform -1 0 4324 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _150_
timestamp -3599
transform -1 0 4232 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _151_
timestamp -3599
transform 1 0 3772 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _152_
timestamp -3599
transform 1 0 4232 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp -3599
transform -1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -3599
transform -1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -3599
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -3599
transform -1 0 2208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp -3599
transform -1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp -3599
transform -1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp -3599
transform -1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp -3599
transform -1 0 3036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp -3599
transform -1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp -3599
transform -1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp -3599
transform -1 0 10028 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp -3599
transform -1 0 9936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp -3599
transform -1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp -3599
transform -1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp -3599
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp -3599
transform -1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp -3599
transform -1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp -3599
transform -1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp -3599
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp -3599
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp -3599
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp -3599
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp -3599
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp -3599
transform -1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp -3599
transform -1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp -3599
transform -1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp -3599
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp -3599
transform -1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp -3599
transform -1 0 10764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp -3599
transform -1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp -3599
transform -1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp -3599
transform -1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp -3599
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform -1 0 8280 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 6716 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 6900 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp -3599
transform 1 0 6716 0 1 4352
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34
timestamp -3599
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp -3599
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp -3599
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70
timestamp -3599
transform 1 0 7544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp -3599
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp -3599
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_8
timestamp -3599
transform 1 0 1840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_16
timestamp -3599
transform 1 0 2576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp -3599
transform 1 0 4600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_64
timestamp -3599
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp -3599
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp -3599
transform 1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp -3599
transform 1 0 6716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp -3599
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_92
timestamp -3599
transform 1 0 9568 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp -3599
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1636964856
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp -3599
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_72
timestamp 1636964856
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp -3599
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1636964856
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_84
timestamp 1636964856
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_10
timestamp 1636964856
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp -3599
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636964856
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp -3599
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp -3599
transform 1 0 2024 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_14
timestamp 1636964856
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1636964856
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1636964856
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp -3599
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp -3599
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_92
timestamp -3599
transform 1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_100
timestamp -3599
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636964856
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_8
timestamp -3599
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_16
timestamp -3599
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1636964856
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_80
timestamp -3599
transform 1 0 8464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp -3599
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp -3599
transform 1 0 10580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_7
timestamp -3599
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_17
timestamp -3599
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp -3599
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636964856
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636964856
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636964856
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp -3599
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp -3599
transform 1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_17
timestamp -3599
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1636964856
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp -3599
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp -3599
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636964856
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636964856
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp -3599
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp -3599
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_100
timestamp -3599
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_6
timestamp -3599
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp -3599
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp -3599
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636964856
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636964856
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636964856
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp -3599
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -3599
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1636964856
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1636964856
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1636964856
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1636964856
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp -3599
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp -3599
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_61
timestamp -3599
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_83
timestamp -3599
transform 1 0 8740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp -3599
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_97
timestamp -3599
transform 1 0 10028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_105
timestamp -3599
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp -3599
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp -3599
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636964856
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636964856
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp -3599
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp -3599
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -3599
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636964856
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_97
timestamp -3599
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_17
timestamp 1636964856
transform 1 0 2668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp -3599
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp -3599
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp -3599
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_72
timestamp -3599
transform 1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_76
timestamp -3599
transform 1 0 8096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_80
timestamp -3599
transform 1 0 8464 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_88
timestamp -3599
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_107
timestamp -3599
transform 1 0 10948 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp -3599
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_18
timestamp -3599
transform 1 0 2760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp -3599
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp -3599
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_50
timestamp 1636964856
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp -3599
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp -3599
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_25
timestamp -3599
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_29
timestamp 1636964856
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp -3599
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_49
timestamp -3599
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp -3599
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp -3599
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp -3599
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_83
timestamp -3599
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp -3599
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_94
timestamp -3599
transform 1 0 9752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform -1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -3599
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -3599
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3599
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -3599
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3599
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -3599
transform 1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -3599
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -3599
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -3599
transform 1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -3599
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -3599
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -3599
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp -3599
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -3599
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -3599
transform 1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp -3599
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp -3599
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp -3599
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp -3599
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp -3599
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp -3599
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp -3599
transform -1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp -3599
transform 1 0 10396 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp -3599
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp -3599
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp -3599
transform -1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp -3599
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp -3599
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_18
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_19
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_20
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_21
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 11316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_22
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_23
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_24
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_25
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_26
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_27
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_28
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_29
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 11316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_30
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_31
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_32
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_33
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_34
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_35
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_40
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_41
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_44
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_45
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_46
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_47
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_48
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_49
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_50
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_51
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_52
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_54
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_55
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_56
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_57
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_58
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_59
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_60
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_62
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_63
timestamp -3599
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_64
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_65
timestamp -3599
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
<< labels >>
flabel metal4 s -2966 -1894 -2346 16038 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 -1894 15386 -1274 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 15418 15386 16038 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14766 -1894 15386 16038 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4868 -1894 5188 16038 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s -2966 6006 15386 6326 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s -2006 -934 -1386 15078 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2006 -934 14426 -314 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2006 14458 14426 15078 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13806 -934 14426 15078 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4208 -1894 4528 16038 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s -2966 5346 15386 5666 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9034 13767 9090 14567 0 FreeSans 224 90 0 0 a_i[0]
port 2 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 a_i[10]
port 3 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 a_i[11]
port 4 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 a_i[12]
port 5 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 a_i[13]
port 6 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 a_i[14]
port 7 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 a_i[15]
port 8 nsew signal input
flabel metal2 s 7746 13767 7802 14567 0 FreeSans 224 90 0 0 a_i[1]
port 9 nsew signal input
flabel metal2 s 6458 13767 6514 14567 0 FreeSans 224 90 0 0 a_i[2]
port 10 nsew signal input
flabel metal3 s 11623 12928 12423 13048 0 FreeSans 480 0 0 0 a_i[3]
port 11 nsew signal input
flabel metal3 s 11623 1368 12423 1488 0 FreeSans 480 0 0 0 a_i[4]
port 12 nsew signal input
flabel metal3 s 11623 2048 12423 2168 0 FreeSans 480 0 0 0 a_i[5]
port 13 nsew signal input
flabel metal3 s 11623 3408 12423 3528 0 FreeSans 480 0 0 0 a_i[6]
port 14 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 a_i[7]
port 15 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 a_i[8]
port 16 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 a_i[9]
port 17 nsew signal input
flabel metal2 s 8390 13767 8446 14567 0 FreeSans 224 90 0 0 b_i[0]
port 18 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 b_i[10]
port 19 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 b_i[11]
port 20 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 b_i[12]
port 21 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 b_i[13]
port 22 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 b_i[14]
port 23 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 b_i[15]
port 24 nsew signal input
flabel metal2 s 7102 13767 7158 14567 0 FreeSans 224 90 0 0 b_i[1]
port 25 nsew signal input
flabel metal3 s 11623 10208 12423 10328 0 FreeSans 480 0 0 0 b_i[2]
port 26 nsew signal input
flabel metal3 s 11623 8168 12423 8288 0 FreeSans 480 0 0 0 b_i[3]
port 27 nsew signal input
flabel metal3 s 11623 5448 12423 5568 0 FreeSans 480 0 0 0 b_i[4]
port 28 nsew signal input
flabel metal3 s 11623 6128 12423 6248 0 FreeSans 480 0 0 0 b_i[5]
port 29 nsew signal input
flabel metal3 s 11623 4088 12423 4208 0 FreeSans 480 0 0 0 b_i[6]
port 30 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 b_i[7]
port 31 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 b_i[8]
port 32 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 b_i[9]
port 33 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 carry_o
port 34 nsew signal output
flabel metal3 s 11623 12248 12423 12368 0 FreeSans 480 0 0 0 clk
port 35 nsew signal input
flabel metal3 s 11623 11568 12423 11688 0 FreeSans 480 0 0 0 sum_o[0]
port 36 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 sum_o[10]
port 37 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 sum_o[11]
port 38 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 sum_o[12]
port 39 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 sum_o[13]
port 40 nsew signal output
flabel metal2 s 5170 13767 5226 14567 0 FreeSans 224 90 0 0 sum_o[14]
port 41 nsew signal output
flabel metal2 s 5814 13767 5870 14567 0 FreeSans 224 90 0 0 sum_o[15]
port 42 nsew signal output
flabel metal3 s 11623 10888 12423 11008 0 FreeSans 480 0 0 0 sum_o[1]
port 43 nsew signal output
flabel metal3 s 11623 9528 12423 9648 0 FreeSans 480 0 0 0 sum_o[2]
port 44 nsew signal output
flabel metal3 s 11623 8848 12423 8968 0 FreeSans 480 0 0 0 sum_o[3]
port 45 nsew signal output
flabel metal3 s 11623 6808 12423 6928 0 FreeSans 480 0 0 0 sum_o[4]
port 46 nsew signal output
flabel metal3 s 11623 7488 12423 7608 0 FreeSans 480 0 0 0 sum_o[5]
port 47 nsew signal output
flabel metal3 s 11623 4768 12423 4888 0 FreeSans 480 0 0 0 sum_o[6]
port 48 nsew signal output
flabel metal3 s 11623 2728 12423 2848 0 FreeSans 480 0 0 0 sum_o[7]
port 49 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 sum_o[8]
port 50 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 sum_o[9]
port 51 nsew signal output
rlabel metal1 6210 11968 6210 11968 0 VGND
rlabel metal1 6210 11424 6210 11424 0 VPWR
rlabel metal2 1886 4964 1886 4964 0 _000_
rlabel metal1 2668 4794 2668 4794 0 _001_
rlabel metal2 2898 4692 2898 4692 0 _002_
rlabel metal1 2116 6766 2116 6766 0 _003_
rlabel metal2 1978 6528 1978 6528 0 _004_
rlabel metal1 2622 6426 2622 6426 0 _005_
rlabel metal1 2760 6834 2760 6834 0 _006_
rlabel metal1 2208 8942 2208 8942 0 _007_
rlabel metal1 2438 8976 2438 8976 0 _008_
rlabel metal2 2254 8330 2254 8330 0 _009_
rlabel metal2 2346 7446 2346 7446 0 _010_
rlabel metal1 2300 10642 2300 10642 0 _011_
rlabel metal1 1840 10574 1840 10574 0 _012_
rlabel metal1 2898 9996 2898 9996 0 _013_
rlabel metal1 2760 10098 2760 10098 0 _014_
rlabel metal1 1932 11118 1932 11118 0 _015_
rlabel metal2 2438 11356 2438 11356 0 _016_
rlabel metal1 3082 11084 3082 11084 0 _017_
rlabel metal1 2254 11186 2254 11186 0 _018_
rlabel metal2 8970 10812 8970 10812 0 _019_
rlabel metal1 7866 10778 7866 10778 0 _020_
rlabel metal1 7958 11186 7958 11186 0 _021_
rlabel metal2 8326 10982 8326 10982 0 _022_
rlabel metal1 7728 10030 7728 10030 0 _023_
rlabel metal2 6854 10268 6854 10268 0 _024_
rlabel metal1 6762 10132 6762 10132 0 _025_
rlabel metal2 7774 9860 7774 9860 0 _026_
rlabel metal2 9154 9452 9154 9452 0 _027_
rlabel metal1 9246 8398 9246 8398 0 _028_
rlabel metal1 9522 9520 9522 9520 0 _029_
rlabel metal2 9246 9180 9246 9180 0 _030_
rlabel metal2 9338 6086 9338 6086 0 _031_
rlabel metal1 9890 6290 9890 6290 0 _032_
rlabel metal2 9338 6596 9338 6596 0 _033_
rlabel metal1 8924 6834 8924 6834 0 _034_
rlabel metal1 8878 5678 8878 5678 0 _035_
rlabel metal2 8694 5440 8694 5440 0 _036_
rlabel metal2 8234 6086 8234 6086 0 _037_
rlabel metal2 8602 5916 8602 5916 0 _038_
rlabel metal1 9798 4114 9798 4114 0 _039_
rlabel metal2 10166 4182 10166 4182 0 _040_
rlabel metal1 9522 4080 9522 4080 0 _041_
rlabel metal2 9430 4794 9430 4794 0 _042_
rlabel metal1 8464 2958 8464 2958 0 _043_
rlabel metal2 8050 2788 8050 2788 0 _044_
rlabel metal2 8786 3332 8786 3332 0 _045_
rlabel metal1 8096 3910 8096 3910 0 _046_
rlabel metal2 5750 3196 5750 3196 0 _047_
rlabel metal1 5520 3162 5520 3162 0 _048_
rlabel metal2 6578 3196 6578 3196 0 _049_
rlabel metal1 6486 2992 6486 2992 0 _050_
rlabel metal2 4094 3332 4094 3332 0 _051_
rlabel metal1 4554 3366 4554 3366 0 _052_
rlabel metal2 4646 3910 4646 3910 0 _053_
rlabel metal1 4002 3468 4002 3468 0 _054_
rlabel metal1 2898 3570 2898 3570 0 _055_
rlabel metal1 1932 4046 1932 4046 0 _056_
rlabel metal1 2438 3468 2438 3468 0 _057_
rlabel metal1 2208 3570 2208 3570 0 _058_
rlabel metal1 2208 5202 2208 5202 0 _059_
rlabel metal2 9062 12828 9062 12828 0 a_i[0]
rlabel metal1 1380 3026 1380 3026 0 a_i[10]
rlabel metal1 1380 4590 1380 4590 0 a_i[11]
rlabel metal1 1380 6290 1380 6290 0 a_i[12]
rlabel via2 1610 9605 1610 9605 0 a_i[13]
rlabel metal1 2208 11730 2208 11730 0 a_i[14]
rlabel metal2 2898 12427 2898 12427 0 a_i[15]
rlabel metal2 7774 12828 7774 12828 0 a_i[1]
rlabel metal2 6486 12828 6486 12828 0 a_i[2]
rlabel metal2 10258 12359 10258 12359 0 a_i[3]
rlabel metal2 10626 1921 10626 1921 0 a_i[4]
rlabel metal2 10350 2261 10350 2261 0 a_i[5]
rlabel via2 10994 3485 10994 3485 0 a_i[6]
rlabel metal2 9062 1520 9062 1520 0 a_i[7]
rlabel metal2 4554 1520 4554 1520 0 a_i[8]
rlabel metal2 3266 1588 3266 1588 0 a_i[9]
rlabel metal2 8418 12828 8418 12828 0 b_i[0]
rlabel metal1 1334 4114 1334 4114 0 b_i[10]
rlabel metal2 1426 5593 1426 5593 0 b_i[11]
rlabel metal3 1004 6868 1004 6868 0 b_i[12]
rlabel metal1 1380 8942 1380 8942 0 b_i[13]
rlabel metal1 1656 10166 1656 10166 0 b_i[14]
rlabel metal1 2438 11730 2438 11730 0 b_i[15]
rlabel metal2 7130 12828 7130 12828 0 b_i[1]
rlabel metal2 10626 10149 10626 10149 0 b_i[2]
rlabel metal2 10626 8143 10626 8143 0 b_i[3]
rlabel metal1 11086 5678 11086 5678 0 b_i[4]
rlabel metal2 10994 6239 10994 6239 0 b_i[5]
rlabel via2 10994 4131 10994 4131 0 b_i[6]
rlabel metal2 7774 1520 7774 1520 0 b_i[7]
rlabel metal2 5842 1520 5842 1520 0 b_i[8]
rlabel metal2 3910 1520 3910 1520 0 b_i[9]
rlabel metal1 1288 11866 1288 11866 0 carry_o
rlabel metal1 9752 7514 9752 7514 0 clk
rlabel metal1 6854 5270 6854 5270 0 clknet_0_clk
rlabel metal1 4094 3570 4094 3570 0 clknet_1_0__leaf_clk
rlabel metal2 4186 8704 4186 8704 0 clknet_1_1__leaf_clk
rlabel metal1 9430 10778 9430 10778 0 fa0.sum_l
rlabel metal1 3112 3094 3112 3094 0 genblk1\[10\].fa0.sum_o
rlabel metal1 3358 5304 3358 5304 0 genblk1\[11\].fa0.sum_o
rlabel metal2 3266 7140 3266 7140 0 genblk1\[12\].fa0.sum_o
rlabel metal1 2714 7990 2714 7990 0 genblk1\[13\].fa0.sum_o
rlabel metal1 3542 10234 3542 10234 0 genblk1\[14\].fa0.sum_o
rlabel metal1 3986 11050 3986 11050 0 genblk1\[15\].fa0.sum_o
rlabel via1 9793 10710 9793 10710 0 genblk1\[1\].fa0.sum_o
rlabel via1 7585 8942 7585 8942 0 genblk1\[2\].fa0.sum_o
rlabel metal1 9690 8874 9690 8874 0 genblk1\[3\].fa0.sum_o
rlabel metal1 9522 6664 9522 6664 0 genblk1\[4\].fa0.sum_o
rlabel metal1 8878 6426 8878 6426 0 genblk1\[5\].fa0.sum_o
rlabel metal2 9890 4386 9890 4386 0 genblk1\[6\].fa0.sum_o
rlabel metal1 9690 3094 9690 3094 0 genblk1\[7\].fa0.sum_o
rlabel metal2 6946 3298 6946 3298 0 genblk1\[8\].fa0.sum_o
rlabel via1 5285 3434 5285 3434 0 genblk1\[9\].fa0.sum_o
rlabel metal2 9338 11322 9338 11322 0 net1
rlabel metal1 9798 9588 9798 9588 0 net10
rlabel metal1 10396 5678 10396 5678 0 net11
rlabel metal1 9246 5202 9246 5202 0 net12
rlabel metal2 10810 3876 10810 3876 0 net13
rlabel metal1 8464 3026 8464 3026 0 net14
rlabel metal2 4738 2822 4738 2822 0 net15
rlabel metal2 3082 2822 3082 2822 0 net16
rlabel metal1 8924 11118 8924 11118 0 net17
rlabel metal2 1702 3706 1702 3706 0 net18
rlabel metal2 1794 5406 1794 5406 0 net19
rlabel metal2 1518 3332 1518 3332 0 net2
rlabel metal1 1932 6290 1932 6290 0 net20
rlabel metal1 1978 8840 1978 8840 0 net21
rlabel metal2 1610 10438 1610 10438 0 net22
rlabel metal1 1794 11764 1794 11764 0 net23
rlabel metal1 7268 11118 7268 11118 0 net24
rlabel metal1 8790 10030 8790 10030 0 net25
rlabel metal2 10074 9044 10074 9044 0 net26
rlabel metal1 10166 5712 10166 5712 0 net27
rlabel via1 8602 5627 8602 5627 0 net28
rlabel metal1 10442 4216 10442 4216 0 net29
rlabel metal2 1610 4998 1610 4998 0 net3
rlabel metal2 8326 2822 8326 2822 0 net30
rlabel metal1 5382 3026 5382 3026 0 net31
rlabel metal1 3542 2380 3542 2380 0 net32
rlabel metal1 1978 11322 1978 11322 0 net33
rlabel metal1 10810 11322 10810 11322 0 net34
rlabel metal2 7222 2652 7222 2652 0 net35
rlabel metal1 5060 2414 5060 2414 0 net36
rlabel metal1 2300 7514 2300 7514 0 net37
rlabel metal1 1702 8500 1702 8500 0 net38
rlabel metal1 5244 10778 5244 10778 0 net39
rlabel metal2 1610 6562 1610 6562 0 net4
rlabel metal2 5658 11526 5658 11526 0 net40
rlabel metal1 10810 10778 10810 10778 0 net41
rlabel metal1 9706 9146 9706 9146 0 net42
rlabel metal2 10994 8636 10994 8636 0 net43
rlabel metal2 10994 7174 10994 7174 0 net44
rlabel metal2 10534 7548 10534 7548 0 net45
rlabel metal2 10994 4998 10994 4998 0 net46
rlabel metal2 10994 2618 10994 2618 0 net47
rlabel metal2 8510 2890 8510 2890 0 net48
rlabel metal1 6486 2414 6486 2414 0 net49
rlabel metal2 1794 9418 1794 9418 0 net5
rlabel metal1 1748 10642 1748 10642 0 net6
rlabel metal1 1978 11696 1978 11696 0 net7
rlabel metal2 7222 11390 7222 11390 0 net8
rlabel metal2 7222 10574 7222 10574 0 net9
rlabel via2 10442 11611 10442 11611 0 sum_o[0]
rlabel metal2 7130 1520 7130 1520 0 sum_o[10]
rlabel metal2 5198 959 5198 959 0 sum_o[11]
rlabel metal3 751 7548 751 7548 0 sum_o[12]
rlabel metal3 1096 8228 1096 8228 0 sum_o[13]
rlabel metal1 5382 11866 5382 11866 0 sum_o[14]
rlabel metal1 5980 11866 5980 11866 0 sum_o[15]
rlabel metal1 11040 11526 11040 11526 0 sum_o[1]
rlabel metal1 11040 9894 11040 9894 0 sum_o[2]
rlabel metal2 10810 8755 10810 8755 0 sum_o[3]
rlabel metal3 11370 6868 11370 6868 0 sum_o[4]
rlabel metal2 10902 7633 10902 7633 0 sum_o[5]
rlabel metal2 10810 4913 10810 4913 0 sum_o[6]
rlabel metal1 10948 2618 10948 2618 0 sum_o[7]
rlabel metal2 8418 1520 8418 1520 0 sum_o[8]
rlabel metal2 6486 1520 6486 1520 0 sum_o[9]
<< properties >>
string FIXED_BBOX 0 0 12423 14567
<< end >>
