* NGSPICE file created from rcAdder.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt rcAdder VGND VPWR a_i[0] a_i[10] a_i[11] a_i[12] a_i[13] a_i[14] a_i[15] a_i[1]
+ a_i[2] a_i[3] a_i[4] a_i[5] a_i[6] a_i[7] a_i[8] a_i[9] b_i[0] b_i[10] b_i[11] b_i[12]
+ b_i[13] b_i[14] b_i[15] b_i[1] b_i[2] b_i[3] b_i[4] b_i[5] b_i[6] b_i[7] b_i[8]
+ b_i[9] carry_o clk sum_o[0] sum_o[10] sum_o[11] sum_o[12] sum_o[13] sum_o[14] sum_o[15]
+ sum_o[1] sum_o[2] sum_o[3] sum_o[4] sum_o[5] sum_o[6] sum_o[7] sum_o[8] sum_o[9]
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_062_ net17 net1 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nand2_1
X_131_ _015_ _016_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ net20 net4 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__or2_1
XANTENNA_input18_A b_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput42 net42 VGND VGND VPWR VPWR sum_o[2] sky130_fd_sc_hd__buf_2
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net23 net7 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nor2_1
X_061_ net24 net8 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__xor2_1
X_113_ _001_ _002_ VGND VGND VPWR VPWR genblk1\[11\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_8_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input30_A b_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput43 net43 VGND VGND VPWR VPWR sum_o[3] sky130_fd_sc_hd__buf_2
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ net24 net8 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and2_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_112_ _055_ _058_ _056_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21bo_1
Xoutput44 net44 VGND VGND VPWR VPWR sum_o[4] sky130_fd_sc_hd__buf_2
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput33 net33 VGND VGND VPWR VPWR carry_o sky130_fd_sc_hd__buf_2
XANTENNA_input23_A b_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_111_ _059_ _000_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nand2_1
Xoutput34 net34 VGND VGND VPWR VPWR sum_o[0] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR sum_o[5] sky130_fd_sc_hd__buf_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input16_A a_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A a_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_110_ net19 net3 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__nand2_1
Xclkload0 clknet_1_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput35 net35 VGND VGND VPWR VPWR sum_o[10] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR sum_o[6] sky130_fd_sc_hd__buf_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput47 net47 VGND VGND VPWR VPWR sum_o[7] sky130_fd_sc_hd__buf_2
Xoutput36 net36 VGND VGND VPWR VPWR sum_o[11] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input21_A b_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_099_ net32 net16 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__or2_1
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput48 net48 VGND VGND VPWR VPWR sum_o[8] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR sum_o[12] sky130_fd_sc_hd__buf_2
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input14_A a_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input6_A a_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ _049_ _050_ VGND VGND VPWR VPWR genblk1\[8\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput49 net49 VGND VGND VPWR VPWR sum_o[9] sky130_fd_sc_hd__buf_2
Xoutput38 net38 VGND VGND VPWR VPWR sum_o[13] sky130_fd_sc_hd__buf_2
XFILLER_15_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ _043_ _046_ _044_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21bo_1
X_149_ clknet_1_1__leaf_clk genblk1\[12\].fa0.sum_o VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
Xoutput39 net39 VGND VGND VPWR VPWR sum_o[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_16_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ _047_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_7_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ clknet_1_0__leaf_clk genblk1\[11\].fa0.sum_o VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_079_ net28 net12 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_A a_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A a_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_095_ net31 net15 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_147_ clknet_1_0__leaf_clk genblk1\[10\].fa0.sum_o VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_078_ _033_ _034_ VGND VGND VPWR VPWR genblk1\[4\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_094_ net31 net15 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or2_1
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_146_ clknet_1_0__leaf_clk genblk1\[9\].fa0.sum_o VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_1
X_077_ _027_ _028_ _029_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a21bo_1
X_129_ net23 net7 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ _045_ _046_ VGND VGND VPWR VPWR genblk1\[7\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
Xinput1 a_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_145_ clknet_1_0__leaf_clk genblk1\[8\].fa0.sum_o VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_1
X_076_ _031_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nand2_1
XANTENNA_input28_A b_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_128_ _013_ _014_ VGND VGND VPWR VPWR genblk1\[14\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input10_A a_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A a_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _039_ _042_ _040_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21bo_1
Xinput2 a_i[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_144_ clknet_1_0__leaf_clk genblk1\[7\].fa0.sum_o VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ net27 net11 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_127_ _007_ _010_ _008_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a21bo_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_091_ _043_ _044_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand2_1
Xinput3 a_i[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_143_ clknet_1_0__leaf_clk genblk1\[6\].fa0.sum_o VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_074_ net27 net11 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__or2_1
XFILLER_7_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_126_ _011_ _012_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ net19 net3 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or2_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ net30 net14 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nand2_1
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 a_i[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_142_ clknet_1_1__leaf_clk genblk1\[5\].fa0.sum_o VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_073_ _027_ _030_ VGND VGND VPWR VPWR genblk1\[3\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_125_ net22 net6 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__nand2_1
XANTENNA_input26_A b_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _057_ _058_ VGND VGND VPWR VPWR genblk1\[10\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 a_i[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_141_ clknet_1_0__leaf_clk genblk1\[4\].fa0.sum_o VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_1
X_072_ _028_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand2_1
XFILLER_7_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_124_ net22 net6 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__or2_1
Xinput30 b_i[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_107_ _051_ _054_ _052_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a21bo_1
XANTENNA_input19_A b_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 a_i[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_140_ clknet_1_1__leaf_clk genblk1\[3\].fa0.sum_o VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_1
X_071_ net26 net10 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput31 b_i[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 b_i[12] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_123_ _009_ _010_ VGND VGND VPWR VPWR genblk1\[13\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_106_ _055_ _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand2_1
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input31_A b_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 a_i[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_070_ net26 net10 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__or2_1
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_122_ _003_ _006_ _004_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 a_i[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 b_i[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput21 b_i[13] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
X_105_ net18 net2 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__nand2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input24_A b_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 a_i[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_121_ _007_ _008_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__nand2_1
Xinput11 a_i[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput22 b_i[14] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
X_104_ net18 net2 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__or2_1
XANTENNA_input17_A b_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A a_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 a_i[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ net21 net5 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nand2_1
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 a_i[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 b_i[15] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_103_ _053_ _054_ VGND VGND VPWR VPWR genblk1\[9\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 b_i[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput13 a_i[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ _047_ _050_ _048_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input22_A b_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 a_i[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 b_i[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
X_101_ _051_ _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nand2_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input15_A a_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input7_A a_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 a_i[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 b_i[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
X_100_ net32 net16 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nand2_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 a_i[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 b_i[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input20_A b_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput17 b_i[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
Xinput28 b_i[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ net30 net14 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__or2_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_input13_A a_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input5_A a_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 b_i[10] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 b_i[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
X_088_ _041_ _042_ VGND VGND VPWR VPWR genblk1\[6\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 b_i[11] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ _035_ _038_ _036_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a21bo_1
X_139_ clknet_1_1__leaf_clk genblk1\[2\].fa0.sum_o VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_086_ _039_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input29_A b_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_069_ _023_ _024_ _025_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21bo_1
X_138_ clknet_1_1__leaf_clk genblk1\[1\].fa0.sum_o VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A a_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input3_A a_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ net29 net13 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_068_ _023_ _026_ VGND VGND VPWR VPWR genblk1\[2\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
X_137_ clknet_1_1__leaf_clk fa0.sum_l VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_12_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_084_ net29 net13 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__or2_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_136_ _022_ _019_ VGND VGND VPWR VPWR fa0.sum_l sky130_fd_sc_hd__and2_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_067_ _024_ _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nand2_1
X_119_ net21 net5 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__or2_1
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_083_ _037_ _038_ VGND VGND VPWR VPWR genblk1\[5\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ clknet_1_1__leaf_clk genblk1\[15\].fa0.sum_o VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
X_066_ net25 net9 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nand2_1
X_135_ net17 net1 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__or2_1
XANTENNA_input27_A b_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_118_ _005_ _006_ VGND VGND VPWR VPWR genblk1\[12\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input1_A a_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _031_ _034_ _032_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a21bo_1
X_151_ clknet_1_1__leaf_clk genblk1\[14\].fa0.sum_o VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ net25 net9 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__or2_1
X_134_ _017_ _018_ VGND VGND VPWR VPWR genblk1\[15\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
X_117_ _059_ _002_ _000_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a21bo_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_081_ _035_ _036_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__nand2_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_150_ clknet_1_1__leaf_clk genblk1\[13\].fa0.sum_o VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_133_ _016_ _018_ _015_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__o21bai_1
X_064_ net17 net1 _021_ _020_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_116_ _003_ _004_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input32_A b_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput40 net40 VGND VGND VPWR VPWR sum_o[15] sky130_fd_sc_hd__buf_2
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_080_ net28 net12 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_132_ _011_ _014_ _012_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21boi_1
X_063_ _021_ _022_ VGND VGND VPWR VPWR genblk1\[1\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ net20 net4 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nand2_1
XANTENNA_input25_A b_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput41 net41 VGND VGND VPWR VPWR sum_o[1] sky130_fd_sc_hd__buf_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

