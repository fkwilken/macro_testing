* NGSPICE file created from rcAdder.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

.subckt rcAdder VGND VPWR a_i[0] a_i[1] a_i[2] a_i[3] b_i[0] b_i[1] b_i[2] b_i[3]
+ carry_o clk sum_o[0] sum_o[1] sum_o[2] sum_o[3]
XTAP_TAPCELL_ROW_8_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR sum_o[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput11 net11 VGND VGND VPWR VPWR sum_o[1] sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput9 net9 VGND VGND VPWR VPWR carry_o sky130_fd_sc_hd__buf_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ clknet_1_1__leaf_clk fa0.sum_l VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
Xoutput12 net12 VGND VGND VPWR VPWR sum_o[2] sky130_fd_sc_hd__buf_2
X_28_ _01_ _02_ VGND VGND VPWR VPWR genblk1\[1\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
Xoutput13 net13 VGND VGND VPWR VPWR sum_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27_ _02_ _11_ VGND VGND VPWR VPWR fa0.sum_l sky130_fd_sc_hd__and2_1
X_26_ net5 net1 VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__or2_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25_ _08_ _10_ VGND VGND VPWR VPWR genblk1\[3\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24_ _08_ _09_ _07_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__o21bai_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23_ _07_ _09_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22_ net8 net4 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_7_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21_ _03_ _04_ _05_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_0_Left_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 a_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_20_ net8 net4 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__and2_1
Xinput2 a_i[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xinput3 a_i[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 a_i[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xinput5 b_i[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_4_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 b_i[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 b_i[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput8 b_i[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19_ _03_ _06_ VGND VGND VPWR VPWR genblk1\[2\].fa0.sum_o sky130_fd_sc_hd__xnor2_1
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18_ _04_ _05_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__nand2_1
X_17_ net7 net3 VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__nand2_1
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16_ net7 net3 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__or2_1
X_15_ net5 net1 _01_ _00_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__a31o_1
X_31_ clknet_1_0__leaf_clk genblk1\[2\].fa0.sum_o VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
X_32_ clknet_1_0__leaf_clk genblk1\[3\].fa0.sum_o VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30_ clknet_1_1__leaf_clk genblk1\[1\].fa0.sum_o VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
X_14_ net5 net1 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ net6 net2 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__and2_1
X_13_ net6 net2 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__xor2_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

