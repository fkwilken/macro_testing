magic
tech sky130A
magscale 1 2
timestamp 1740619358
<< viali >>
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3985 6681 4019 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 5273 6613 5307 6647
rect 1593 6273 1627 6307
rect 2237 6273 2271 6307
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 5365 6273 5399 6307
rect 5733 6273 5767 6307
rect 1685 6205 1719 6239
rect 2421 6205 2455 6239
rect 5549 6137 5583 6171
rect 1961 6069 1995 6103
rect 2053 6069 2087 6103
rect 2605 6069 2639 6103
rect 5181 6069 5215 6103
rect 1593 5865 1627 5899
rect 5733 5865 5767 5899
rect 2053 5729 2087 5763
rect 2237 5729 2271 5763
rect 2329 5729 2363 5763
rect 2697 5729 2731 5763
rect 3249 5729 3283 5763
rect 4353 5729 4387 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 3433 5661 3467 5695
rect 4598 5593 4632 5627
rect 1869 5525 1903 5559
rect 2513 5525 2547 5559
rect 3157 5525 3191 5559
rect 3617 5525 3651 5559
rect 2881 5321 2915 5355
rect 5733 5321 5767 5355
rect 2513 5253 2547 5287
rect 2697 5253 2731 5287
rect 4598 5253 4632 5287
rect 1409 5185 1443 5219
rect 4353 5185 4387 5219
rect 1593 4981 1627 5015
rect 4261 4777 4295 4811
rect 1869 4641 1903 4675
rect 1409 4573 1443 4607
rect 1777 4573 1811 4607
rect 1961 4573 1995 4607
rect 2329 4573 2363 4607
rect 2513 4573 2547 4607
rect 5733 4573 5767 4607
rect 1593 4437 1627 4471
rect 2513 4437 2547 4471
rect 1593 4165 1627 4199
rect 1777 4165 1811 4199
rect 2053 4097 2087 4131
rect 2421 4097 2455 4131
rect 2513 4097 2547 4131
rect 2789 4097 2823 4131
rect 4609 4097 4643 4131
rect 2881 4029 2915 4063
rect 4353 4029 4387 4063
rect 1961 3961 1995 3995
rect 3157 3961 3191 3995
rect 2237 3893 2271 3927
rect 5733 3893 5767 3927
rect 2605 3553 2639 3587
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 2053 3485 2087 3519
rect 2237 3485 2271 3519
rect 2697 3485 2731 3519
rect 4353 3485 4387 3519
rect 4598 3417 4632 3451
rect 1501 3349 1535 3383
rect 1961 3349 1995 3383
rect 3065 3349 3099 3383
rect 5733 3349 5767 3383
rect 1777 3145 1811 3179
rect 2329 3145 2363 3179
rect 5181 3145 5215 3179
rect 5549 3145 5583 3179
rect 2605 3077 2639 3111
rect 1409 3009 1443 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2421 3009 2455 3043
rect 2513 3009 2547 3043
rect 2697 3009 2731 3043
rect 5365 3009 5399 3043
rect 5733 3009 5767 3043
rect 2145 2941 2179 2975
rect 1593 2873 1627 2907
rect 1593 2601 1627 2635
rect 5273 2601 5307 2635
rect 1409 2397 1443 2431
rect 3985 2397 4019 2431
<< metal1 >>
rect 1104 7098 6072 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 6072 7098
rect 1104 7024 6072 7046
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 992 6752 1409 6780
rect 992 6740 998 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1397 6743 1455 6749
rect 1504 6752 1685 6780
rect 842 6672 848 6724
rect 900 6712 906 6724
rect 1504 6712 1532 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 2222 6712 2228 6724
rect 900 6684 1532 6712
rect 1596 6684 2228 6712
rect 900 6672 906 6684
rect 1596 6653 1624 6684
rect 2222 6672 2228 6684
rect 2280 6712 2286 6724
rect 2498 6712 2504 6724
rect 2280 6684 2504 6712
rect 2280 6672 2286 6684
rect 2498 6672 2504 6684
rect 2556 6672 2562 6724
rect 3970 6672 3976 6724
rect 4028 6672 4034 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 4396 6616 5273 6644
rect 4396 6604 4402 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 1104 6554 6072 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 6072 6554
rect 1104 6480 6072 6502
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 1728 6344 2268 6372
rect 1728 6332 1734 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1854 6304 1860 6316
rect 1627 6276 1860 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1854 6264 1860 6276
rect 1912 6304 1918 6316
rect 2240 6313 2268 6344
rect 2225 6307 2283 6313
rect 1912 6276 1992 6304
rect 1912 6264 1918 6276
rect 1670 6196 1676 6248
rect 1728 6196 1734 6248
rect 1964 6236 1992 6276
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5626 6304 5632 6316
rect 5399 6276 5632 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 2409 6239 2467 6245
rect 2409 6236 2421 6239
rect 1964 6208 2421 6236
rect 2409 6205 2421 6208
rect 2455 6205 2467 6239
rect 2409 6199 2467 6205
rect 5534 6128 5540 6180
rect 5592 6128 5598 6180
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 2038 6060 2044 6112
rect 2096 6060 2102 6112
rect 2593 6103 2651 6109
rect 2593 6069 2605 6103
rect 2639 6100 2651 6103
rect 2682 6100 2688 6112
rect 2639 6072 2688 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5902 6100 5908 6112
rect 5215 6072 5908 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 1104 6010 6072 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 6072 6010
rect 1104 5936 6072 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1670 5896 1676 5908
rect 1627 5868 1676 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 5718 5856 5724 5908
rect 5776 5856 5782 5908
rect 1946 5788 1952 5840
rect 2004 5828 2010 5840
rect 2004 5800 2360 5828
rect 2004 5788 2010 5800
rect 2038 5720 2044 5772
rect 2096 5720 2102 5772
rect 2222 5720 2228 5772
rect 2280 5720 2286 5772
rect 2332 5769 2360 5800
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 900 5664 1409 5692
rect 900 5652 906 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2332 5692 2360 5723
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3237 5763 3295 5769
rect 3237 5760 3249 5763
rect 2740 5732 3249 5760
rect 2740 5720 2746 5732
rect 3237 5729 3249 5732
rect 3283 5729 3295 5763
rect 3237 5723 3295 5729
rect 4338 5720 4344 5772
rect 4396 5720 4402 5772
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2332 5664 2789 5692
rect 2133 5655 2191 5661
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2148 5624 2176 5655
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 2682 5624 2688 5636
rect 2148 5596 2688 5624
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 2148 5556 2176 5596
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 4586 5627 4644 5633
rect 4586 5624 4598 5627
rect 3160 5596 4598 5624
rect 1903 5528 2176 5556
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 3160 5565 3188 5596
rect 4586 5593 4598 5596
rect 4632 5593 4644 5627
rect 4586 5587 4644 5593
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2280 5528 2513 5556
rect 2280 5516 2286 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3605 5559 3663 5565
rect 3605 5525 3617 5559
rect 3651 5556 3663 5559
rect 4430 5556 4436 5568
rect 3651 5528 4436 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 1104 5466 6072 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 6072 5466
rect 1104 5392 6072 5414
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3418 5352 3424 5364
rect 2915 5324 3424 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5684 5324 5733 5352
rect 5684 5312 5690 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 2314 5244 2320 5296
rect 2372 5284 2378 5296
rect 2501 5287 2559 5293
rect 2501 5284 2513 5287
rect 2372 5256 2513 5284
rect 2372 5244 2378 5256
rect 2501 5253 2513 5256
rect 2547 5253 2559 5287
rect 2501 5247 2559 5253
rect 2682 5244 2688 5296
rect 2740 5244 2746 5296
rect 4430 5244 4436 5296
rect 4488 5284 4494 5296
rect 4586 5287 4644 5293
rect 4586 5284 4598 5287
rect 4488 5256 4598 5284
rect 4488 5244 4494 5256
rect 4586 5253 4598 5256
rect 4632 5253 4644 5287
rect 4586 5247 4644 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 1946 5012 1952 5024
rect 1627 4984 1952 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 1104 4922 6072 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 6072 4922
rect 1104 4848 6072 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4028 4780 4261 4808
rect 4028 4768 4034 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 2038 4672 2044 4684
rect 1903 4644 2044 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2038 4632 2044 4644
rect 2096 4672 2102 4684
rect 2096 4644 2360 4672
rect 2096 4632 2102 4644
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1397 4567 1455 4573
rect 1596 4576 1777 4604
rect 1596 4480 1624 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 1946 4564 1952 4616
rect 2004 4564 2010 4616
rect 2332 4613 2360 4644
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2498 4564 2504 4616
rect 2556 4564 2562 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 2501 4471 2559 4477
rect 2501 4437 2513 4471
rect 2547 4468 2559 4471
rect 2866 4468 2872 4480
rect 2547 4440 2872 4468
rect 2547 4437 2559 4440
rect 2501 4431 2559 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 1104 4378 6072 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 6072 4378
rect 1104 4304 6072 4326
rect 1578 4156 1584 4208
rect 1636 4156 1642 4208
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4196 1823 4199
rect 1946 4196 1952 4208
rect 1811 4168 1952 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 2038 4088 2044 4140
rect 2096 4088 2102 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 2280 4100 2421 4128
rect 2280 4088 2286 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2424 4060 2452 4091
rect 2498 4088 2504 4140
rect 2556 4088 2562 4140
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 4597 4131 4655 4137
rect 4597 4128 4609 4131
rect 2777 4091 2835 4097
rect 3804 4100 4609 4128
rect 2792 4060 2820 4091
rect 2424 4032 2820 4060
rect 2866 4020 2872 4072
rect 2924 4020 2930 4072
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2498 3992 2504 4004
rect 1995 3964 2504 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3804 3992 3832 4100
rect 4597 4097 4609 4100
rect 4643 4097 4655 4131
rect 4597 4091 4655 4097
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 3191 3964 3832 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 1104 3834 6072 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 6072 3834
rect 1104 3760 6072 3782
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2593 3587 2651 3593
rect 2593 3584 2605 3587
rect 2372 3556 2605 3584
rect 2372 3544 2378 3556
rect 2593 3553 2605 3556
rect 2639 3553 2651 3587
rect 2593 3547 2651 3553
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1688 3448 1716 3479
rect 1762 3476 1768 3528
rect 1820 3476 1826 3528
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2056 3448 2084 3479
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2280 3488 2697 3516
rect 2280 3476 2286 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 4338 3476 4344 3528
rect 4396 3476 4402 3528
rect 2406 3448 2412 3460
rect 1688 3420 1992 3448
rect 2056 3420 2412 3448
rect 842 3340 848 3392
rect 900 3380 906 3392
rect 1964 3389 1992 3420
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 4586 3451 4644 3457
rect 4586 3448 4598 3451
rect 3068 3420 4598 3448
rect 3068 3389 3096 3420
rect 4586 3417 4598 3420
rect 4632 3417 4644 3451
rect 4586 3411 4644 3417
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 900 3352 1501 3380
rect 900 3340 906 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 1489 3343 1547 3349
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3349 2007 3383
rect 1949 3343 2007 3349
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 5721 3383 5779 3389
rect 5721 3349 5733 3383
rect 5767 3380 5779 3383
rect 5767 3352 6132 3380
rect 5767 3349 5779 3352
rect 5721 3343 5779 3349
rect 1104 3290 6072 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 6072 3290
rect 1104 3216 6072 3238
rect 1762 3136 1768 3188
rect 1820 3136 1826 3188
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 1780 3108 1808 3136
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 1780 3080 2268 3108
rect 842 3000 848 3052
rect 900 3040 906 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 900 3012 1409 3040
rect 900 3000 906 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2240 3049 2268 3080
rect 2424 3080 2605 3108
rect 2424 3052 2452 3080
rect 2593 3077 2605 3080
rect 2639 3077 2651 3111
rect 6104 3108 6132 3352
rect 2593 3071 2651 3077
rect 5368 3080 6132 3108
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 5368 3049 5396 3080
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2700 2972 2728 3003
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 2179 2944 2728 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 2148 2904 2176 2935
rect 1627 2876 2176 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 2498 2836 2504 2848
rect 2004 2808 2504 2836
rect 2004 2796 2010 2808
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 1104 2746 6072 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 6072 2746
rect 1104 2672 6072 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 1946 2632 1952 2644
rect 1627 2604 1952 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 4396 2604 5273 2632
rect 4396 2592 4402 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 1104 2202 6072 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 6072 2202
rect 1104 2128 6072 2150
<< via1 >>
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 940 6740 992 6792
rect 848 6672 900 6724
rect 2228 6672 2280 6724
rect 2504 6672 2556 6724
rect 3976 6715 4028 6724
rect 3976 6681 3985 6715
rect 3985 6681 4019 6715
rect 4019 6681 4028 6715
rect 3976 6672 4028 6681
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 4344 6604 4396 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 1676 6332 1728 6384
rect 1860 6264 1912 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 5632 6264 5684 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5540 6171 5592 6180
rect 5540 6137 5549 6171
rect 5549 6137 5583 6171
rect 5583 6137 5592 6171
rect 5540 6128 5592 6137
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 2688 6060 2740 6112
rect 5908 6060 5960 6112
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 1676 5856 1728 5908
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 1952 5788 2004 5840
rect 2044 5763 2096 5772
rect 2044 5729 2053 5763
rect 2053 5729 2087 5763
rect 2087 5729 2096 5763
rect 2044 5720 2096 5729
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 848 5652 900 5704
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 2688 5584 2740 5636
rect 2228 5516 2280 5568
rect 4436 5516 4488 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 3424 5312 3476 5364
rect 5632 5312 5684 5364
rect 2320 5244 2372 5296
rect 2688 5287 2740 5296
rect 2688 5253 2697 5287
rect 2697 5253 2731 5287
rect 2731 5253 2740 5287
rect 2688 5244 2740 5253
rect 4436 5244 4488 5296
rect 848 5176 900 5228
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 1952 4972 2004 5024
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 3976 4768 4028 4820
rect 2044 4632 2096 4684
rect 848 4564 900 4616
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2872 4428 2924 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 1584 4199 1636 4208
rect 1584 4165 1593 4199
rect 1593 4165 1627 4199
rect 1627 4165 1636 4199
rect 1584 4156 1636 4165
rect 1952 4156 2004 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2228 4088 2280 4140
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 2504 3952 2556 4004
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 4344 4020 4396 4029
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 2320 3544 2372 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 848 3340 900 3392
rect 2412 3408 2464 3460
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 848 3000 900 3052
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 1952 2796 2004 2848
rect 2504 2796 2556 2848
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 1952 2592 2004 2644
rect 4344 2592 4396 2644
rect 848 2388 900 2440
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
<< metal2 >>
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 952 6798 980 7511
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 940 6792 992 6798
rect 846 6760 902 6769
rect 940 6734 992 6740
rect 846 6695 848 6704
rect 900 6695 902 6704
rect 2228 6724 2280 6730
rect 848 6666 900 6672
rect 2228 6666 2280 6672
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 1688 6254 1716 6326
rect 1872 6322 1900 6598
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 860 5710 888 6015
rect 1688 5914 1716 6190
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1964 5846 1992 6054
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 2056 5778 2084 6054
rect 2240 5778 2268 6666
rect 2516 6322 2544 6666
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 6202 2728 6258
rect 2700 6174 2820 6202
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 2700 5778 2728 6054
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2240 5658 2268 5714
rect 2792 5658 2820 6174
rect 1688 5545 1716 5646
rect 2240 5630 2360 5658
rect 2700 5642 2820 5658
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 2228 5568 2280 5574
rect 1674 5536 1730 5545
rect 2228 5510 2280 5516
rect 1674 5471 1730 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 1952 5024 2004 5030
rect 846 4992 902 5001
rect 1952 4966 2004 4972
rect 846 4927 902 4936
rect 1964 4622 1992 4966
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 860 4321 888 4558
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 1596 4214 1624 4422
rect 1964 4214 1992 4558
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2056 4146 2084 4626
rect 2240 4146 2268 5510
rect 2332 5302 2360 5630
rect 2688 5636 2820 5642
rect 2740 5630 2820 5636
rect 2688 5578 2740 5584
rect 2700 5302 2728 5578
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3436 5370 3464 5646
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 3988 4826 4016 6666
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 5778 4384 6598
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5538 6216 5594 6225
rect 5538 6151 5540 6160
rect 5592 6151 5594 6160
rect 5540 6122 5592 6128
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5234 4384 5714
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5302 4476 5510
rect 5644 5370 5672 6258
rect 5736 5914 5764 6258
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5920 5545 5948 6054
rect 5906 5536 5962 5545
rect 5906 5471 5962 5480
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 5722 4856 5778 4865
rect 3976 4820 4028 4826
rect 5722 4791 5778 4800
rect 3976 4762 4028 4768
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2516 4146 2544 4558
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 4010 2544 4082
rect 2884 4078 2912 4422
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3534 2268 3878
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 848 3392 900 3398
rect 846 3360 848 3369
rect 900 3360 902 3369
rect 846 3295 902 3304
rect 1780 3194 1808 3470
rect 2332 3194 2360 3538
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2424 3058 2452 3402
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 848 3052 900 3058
rect 848 2994 900 3000
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 860 2961 888 2994
rect 846 2952 902 2961
rect 846 2887 902 2896
rect 1964 2854 1992 2994
rect 2516 2854 2544 2994
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 1964 2650 1992 2790
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 3988 2446 4016 4762
rect 5736 4622 5764 4791
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3534 4384 4014
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 5170 3496 5226 3505
rect 4356 2650 4384 3470
rect 5170 3431 5226 3440
rect 5184 3194 5212 3431
rect 5552 3194 5580 4111
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5736 3058 5764 3878
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 860 2281 888 2382
rect 846 2272 902 2281
rect 846 2207 902 2216
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
<< via2 >>
rect 938 7520 994 7576
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 846 6724 902 6760
rect 846 6704 848 6724
rect 848 6704 900 6724
rect 900 6704 902 6724
rect 846 6024 902 6080
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 1674 5480 1730 5536
rect 846 4936 902 4992
rect 846 4256 902 4312
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 5538 6180 5594 6216
rect 5538 6160 5540 6180
rect 5540 6160 5592 6180
rect 5592 6160 5594 6180
rect 5906 5480 5962 5536
rect 5722 4800 5778 4856
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 846 3340 848 3360
rect 848 3340 900 3360
rect 900 3340 902 3360
rect 846 3304 902 3340
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 846 2896 902 2952
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 5538 4120 5594 4176
rect 5170 3440 5226 3496
rect 846 2216 902 2272
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
<< metal3 >>
rect 0 7578 800 7608
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 0 6898 800 6928
rect 0 6808 858 6898
rect 798 6765 858 6808
rect 798 6760 907 6765
rect 798 6704 846 6760
rect 902 6704 907 6760
rect 798 6702 907 6704
rect 841 6699 907 6702
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 0 6218 800 6248
rect 5533 6218 5599 6221
rect 6385 6218 7185 6248
rect 0 6128 858 6218
rect 5533 6216 7185 6218
rect 5533 6160 5538 6216
rect 5594 6160 7185 6216
rect 5533 6158 7185 6160
rect 5533 6155 5599 6158
rect 6385 6128 7185 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 0 5538 800 5568
rect 1669 5538 1735 5541
rect 0 5536 1735 5538
rect 0 5480 1674 5536
rect 1730 5480 1735 5536
rect 0 5478 1735 5480
rect 0 5448 800 5478
rect 1669 5475 1735 5478
rect 5901 5538 5967 5541
rect 6385 5538 7185 5568
rect 5901 5536 7185 5538
rect 5901 5480 5906 5536
rect 5962 5480 7185 5536
rect 5901 5478 7185 5480
rect 5901 5475 5967 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 6385 5448 7185 5478
rect 3006 5407 3322 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 2346 4928 2662 4929
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 5717 4858 5783 4861
rect 6385 4858 7185 4888
rect 5717 4856 7185 4858
rect 5717 4800 5722 4856
rect 5778 4800 7185 4856
rect 5717 4798 7185 4800
rect 0 4768 800 4798
rect 5717 4795 5783 4798
rect 6385 4768 7185 4798
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 5533 4178 5599 4181
rect 6385 4178 7185 4208
rect 5533 4176 7185 4178
rect 5533 4120 5538 4176
rect 5594 4120 7185 4176
rect 5533 4118 7185 4120
rect 0 4088 800 4118
rect 5533 4115 5599 4118
rect 6385 4088 7185 4118
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 0 3498 800 3528
rect 5165 3498 5231 3501
rect 6385 3498 7185 3528
rect 0 3408 858 3498
rect 5165 3496 7185 3498
rect 5165 3440 5170 3496
rect 5226 3440 7185 3496
rect 5165 3438 7185 3440
rect 5165 3435 5231 3438
rect 6385 3408 7185 3438
rect 798 3365 858 3408
rect 798 3360 907 3365
rect 798 3304 846 3360
rect 902 3304 907 3360
rect 798 3302 907 3304
rect 841 3299 907 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 0 2728 800 2758
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 2346 2687 2662 2688
rect 841 2274 907 2277
rect 798 2272 907 2274
rect 798 2216 846 2272
rect 902 2216 907 2272
rect 798 2211 907 2216
rect 798 2168 858 2211
rect 0 2078 858 2168
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 0 2048 800 2078
<< via3 >>
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
<< metal4 >>
rect 2344 7104 2664 7120
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 2752 2664 3776
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 2128 2664 2688
rect 3004 6560 3324 7120
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 2128 3324 2144
use sky130_fd_sc_hd__and2_1  _12_
timestamp -3599
transform -1 0 2484 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _13_
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _14_
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _15_
timestamp -3599
transform -1 0 2576 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _16_
timestamp -3599
transform 1 0 1564 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _17_
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _18_
timestamp -3599
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp -3599
transform 1 0 2576 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _20_
timestamp -3599
transform -1 0 2208 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _21_
timestamp -3599
transform 1 0 2024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _22_
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _23_
timestamp -3599
transform -1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _24_
timestamp -3599
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _25_
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _26_
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _27_
timestamp -3599
transform 1 0 3220 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _28_
timestamp -3599
transform 1 0 2576 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp -3599
transform 1 0 4324 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp -3599
transform 1 0 4324 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform -1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 3956 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 3956 0 1 6528
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6
timestamp 1636964856
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp -3599
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1636964856
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1636964856
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp -3599
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp -3599
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1636964856
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_10
timestamp -3599
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_16
timestamp 1636964856
transform 1 0 2576 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_14
timestamp -3599
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1636964856
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_32
timestamp -3599
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_18
timestamp 1636964856
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_30
timestamp 1636964856
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_9
timestamp 1636964856
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -3599
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -3599
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3599
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3599
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -3599
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -3599
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform -1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform -1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform -1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_9
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_10
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_11
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_12
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_13
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_14
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 6072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_15
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_16
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_17
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_18
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_19
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_20
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_21
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_22
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
<< labels >>
flabel metal4 s 3004 2128 3324 7120 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2344 2128 2664 7120 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 a_i[0]
port 2 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 a_i[1]
port 3 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 a_i[2]
port 4 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 a_i[3]
port 5 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 b_i[0]
port 6 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 b_i[1]
port 7 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 b_i[2]
port 8 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 b_i[3]
port 9 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 carry_o
port 10 nsew signal output
flabel metal3 s 6385 4768 7185 4888 0 FreeSans 480 0 0 0 clk
port 11 nsew signal input
flabel metal3 s 6385 5448 7185 5568 0 FreeSans 480 0 0 0 sum_o[0]
port 12 nsew signal output
flabel metal3 s 6385 6128 7185 6248 0 FreeSans 480 0 0 0 sum_o[1]
port 13 nsew signal output
flabel metal3 s 6385 4088 7185 4208 0 FreeSans 480 0 0 0 sum_o[2]
port 14 nsew signal output
flabel metal3 s 6385 3408 7185 3528 0 FreeSans 480 0 0 0 sum_o[3]
port 15 nsew signal output
rlabel metal1 3588 6528 3588 6528 0 VGND
rlabel metal1 3588 7072 3588 7072 0 VPWR
rlabel metal2 2070 5916 2070 5916 0 _00_
rlabel metal1 2346 5780 2346 5780 0 _01_
rlabel metal2 2714 5916 2714 5916 0 _02_
rlabel metal1 2346 4114 2346 4114 0 _03_
rlabel metal2 2530 4046 2530 4046 0 _04_
rlabel metal1 2346 4624 2346 4624 0 _05_
rlabel metal2 2898 4250 2898 4250 0 _06_
rlabel metal2 1794 3332 1794 3332 0 _07_
rlabel metal2 2254 3706 2254 3706 0 _08_
rlabel metal2 2438 3230 2438 3230 0 _09_
rlabel metal2 2346 3366 2346 3366 0 _10_
rlabel metal1 3174 5338 3174 5338 0 _11_
rlabel metal1 1196 6766 1196 6766 0 a_i[0]
rlabel metal3 751 6188 751 6188 0 a_i[1]
rlabel metal3 751 4148 751 4148 0 a_i[2]
rlabel metal3 751 2108 751 2108 0 a_i[3]
rlabel metal3 1188 5508 1188 5508 0 b_i[0]
rlabel metal3 751 6868 751 6868 0 b_i[1]
rlabel metal3 751 4828 751 4828 0 b_i[2]
rlabel metal3 751 2788 751 2788 0 b_i[3]
rlabel metal3 751 3468 751 3468 0 carry_o
rlabel metal2 5750 4709 5750 4709 0 clk
rlabel metal1 4140 4794 4140 4794 0 clknet_0_clk
rlabel metal2 4370 3060 4370 3060 0 clknet_1_0__leaf_clk
rlabel metal2 4370 6188 4370 6188 0 clknet_1_1__leaf_clk
rlabel metal1 4538 5270 4538 5270 0 fa0.sum_l
rlabel metal1 3894 5610 3894 5610 0 genblk1\[1\].fa0.sum_o
rlabel metal1 3496 3978 3496 3978 0 genblk1\[2\].fa0.sum_o
rlabel metal1 3848 3434 3848 3434 0 genblk1\[3\].fa0.sum_o
rlabel metal2 2530 6494 2530 6494 0 net1
rlabel metal1 5704 5338 5704 5338 0 net10
rlabel metal2 5750 6086 5750 6086 0 net11
rlabel metal2 5750 3468 5750 3468 0 net12
rlabel metal1 5382 3060 5382 3060 0 net13
rlabel metal2 1702 6052 1702 6052 0 net2
rlabel metal1 1702 4590 1702 4590 0 net3
rlabel via1 1978 2822 1978 2822 0 net4
rlabel metal2 2714 5457 2714 5457 0 net5
rlabel metal1 1794 6290 1794 6290 0 net6
rlabel metal2 1978 4794 1978 4794 0 net7
rlabel metal1 2162 2924 2162 2924 0 net8
rlabel metal1 1702 3468 1702 3468 0 net9
rlabel metal1 5566 6086 5566 6086 0 sum_o[0]
rlabel via2 5566 6171 5566 6171 0 sum_o[1]
rlabel metal2 5566 3655 5566 3655 0 sum_o[2]
rlabel metal2 5198 3315 5198 3315 0 sum_o[3]
<< properties >>
string FIXED_BBOX 0 0 7185 9329
<< end >>
