VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rcAdder
  CLASS BLOCK ;
  FOREIGN rcAdder ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.925 BY 46.645 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 35.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 35.600 ;
    END
  END VPWR
  PIN a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a_i[0]
  PIN a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END a_i[1]
  PIN a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a_i[2]
  PIN a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END a_i[3]
  PIN b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b_i[0]
  PIN b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b_i[1]
  PIN b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END b_i[2]
  PIN b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END b_i[3]
  PIN carry_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END carry_o
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 31.925 23.840 35.925 24.440 ;
    END
  END clk
  PIN sum_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 31.925 27.240 35.925 27.840 ;
    END
  END sum_o[0]
  PIN sum_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 31.925 30.640 35.925 31.240 ;
    END
  END sum_o[1]
  PIN sum_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 31.925 20.440 35.925 21.040 ;
    END
  END sum_o[2]
  PIN sum_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 31.925 17.040 35.925 17.640 ;
    END
  END sum_o[3]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 30.550 35.550 ;
      LAYER li1 ;
        RECT 5.520 10.795 30.360 35.445 ;
      LAYER met1 ;
        RECT 4.210 10.640 30.660 35.600 ;
      LAYER met2 ;
        RECT 4.230 10.695 29.810 37.925 ;
      LAYER met3 ;
        RECT 4.400 37.040 31.925 37.905 ;
        RECT 3.990 35.040 31.925 37.040 ;
        RECT 4.400 33.640 31.925 35.040 ;
        RECT 3.990 31.640 31.925 33.640 ;
        RECT 4.400 30.240 31.525 31.640 ;
        RECT 3.990 28.240 31.925 30.240 ;
        RECT 4.400 26.840 31.525 28.240 ;
        RECT 3.990 24.840 31.925 26.840 ;
        RECT 4.400 23.440 31.525 24.840 ;
        RECT 3.990 21.440 31.925 23.440 ;
        RECT 4.400 20.040 31.525 21.440 ;
        RECT 3.990 18.040 31.925 20.040 ;
        RECT 4.400 16.640 31.525 18.040 ;
        RECT 3.990 14.640 31.925 16.640 ;
        RECT 4.400 13.240 31.925 14.640 ;
        RECT 3.990 11.240 31.925 13.240 ;
        RECT 4.400 10.390 31.925 11.240 ;
  END
END rcAdder
END LIBRARY

